/*
	Copyright 2020 Mohamed Shalan (mshalan@aucegypt.edu)
	
	Licensed under the Apache License, Version 2.0 (the "License"); 
	you may not use this file except in compliance with the License. 
	You may obtain a copy of the License at:
	http://www.apache.org/licenses/LICENSE-2.0
	Unless required by applicable law or agreed to in writing, software 
	distributed under the License is distributed on an "AS IS" BASIS, 
	WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
	See the License for the specific language governing permissions and 
	limitations under the License.
*/

`timescale              1ns/1ps
`default_nettype        none

/* 
    Clock and Reset Manager 
     - Internal RC Oscillator (2mhz, 8mhz, 16mhz)
     - Clock Multiplexor
     - Clock divider (/2, /4, /8 and /16)
*/
module MS_CLK_RST(
    `ifdef GL 
        input   wire    vccd1,
        input   wire    vssd1,
    `endif // GL
    input   wire        xclk,           // External clock source 
    input   wire        xrst_n,         // external reset
    input   wire        por_n,          // Power-on-Reset
    input   wire        dll_en,         // Enable DLL
    input   wire [4:0]  dll_div,        // DLL feedback division ratio
    input   wire        dll_dco,        // Run in DCO mode
    input   wire [25:0] dll_ext_trim,   // External trim for DCO mode
    input   wire        sel_mux0,       // CLKMUX0 selection - 0: ROSC 16MHz    1: ROSC 2MHz
    input   wire        sel_mux1,       // CLKMUX1 selection - 0: dll_clk       1: XCLK
    input   wire        sel_mux2,       // CLKMUX2 selection - 0: ROSC 16 or 2  1: XCLK or dll
    input   wire        sel_mux3,       // CLKMUX3 selection - 0: CLKMUX2 div   1: CLKMUX2 output
    input   wire        sel_mux4,       // CLKMUX4 selection - 0: ROSC 8MHz     1: CLKMUX3 output
    input   wire [1:0]  rosc_en,        // ROSC Enable: 8MHz is generated by default; bit 0: 2MHz enable, bit 1: 16MHz enable
    input   wire [3:0]  rosc_trim,      // ROSC trim: bit 1-0: 2MHz trim, bit 3-2: 16MHz trim
    input   wire [1:0]  clk_div,        // Clock divider for the output of CLKMUX2: 2, 4, 8 and 16

    output  wire        clk,            // system clock
    output  wire        clk_div_2,          // system clock divided by 2
    output  wire        rst_n           // system reset
);

    wire clk_2mhz, clk_8mhz, clk_16mhz;
    rosc ROSC(
    `ifdef PnR
        VGND(VGND),
        VNB(VNB),
        VPB(VPB),
        VPWR(VPWR),
    `endif // PnR
        .en_2mhz(rosc_en[0]),
        .en_16mhz(rosc_en[1]),
        .trim_2mhz(rosc_trim[1:0]),
        .trim_16mhz(rosc_trim[3:2]),
        .clk_2mhz(clk_2mhz),
        .clk_8mhz(clk_8mhz),
        .clk_16mhz(clk_16mhz)
    );

    // internal reset logic
    wire    irst_n;

    assign irst_n = xrst_n & por_n;

    // Reset Synchonizer
    rst_sync RST_SYNC (
	    .clk(clk_8mhz),
	    .rst_n(irst_n),
	    .srst_n(rst_n)
    );

    wire    clk_mux0;
    clkmux_2x1 CLKMUX0 (
        .rst_n(rst_n),
        .clk0(clk_16mhz), 
        .clk1(clk_2mhz), 
        .sel(sel_mux0),
        .clko(clk_mux0)
    );

    /* Internally generated clock */
    wire dll_clk, dll_clk90;
    digital_locked_loop dll (
        .resetb(rst_n),
        .enable(dll_en),
        .osc(xclk),
        .clockp({dll_clk, dll_clk90}),
        .div(dll_div),
        .dco(dll_dco),
        .ext_trim(dll_ext_trim)
    );

    wire    clk_mux1;
    clkmux_2x1 CLKMUX1 (
        .rst_n(rst_n),
        .clk0(dll_clk), 
        .clk1(xclk), 
        .sel(sel_mux1),
        .clko(clk_mux1)
    );
        
    wire    clk_mux2;
    clkmux_2x1 CLKMUX2 (
        .rst_n(rst_n),
        .clk0(clk_mux0), 
        .clk1(clk_mux1), 
        .sel(sel_mux2),
        .clko(clk_mux2)
    );

    // Clock Divider
    reg [3:0]   clkdiv = 0;
    always@(posedge clk_mux2)
        clkdiv <= clkdiv + 1'b1;

    wire    clk_2   = clkdiv[0];
    wire    clk_4   = clkdiv[1];
    wire    clk_8   = clkdiv[2];
    wire    clk_16  = clkdiv[3];
    
    wire    clk_mux2_div;
    clkmux_4x1 CLKMUX (
        .rst_n(rst_n),
        .clk0(clk_2), 
        .clk1(clk_4), 
        .clk2(clk_8),
        .clk3(clk_16),
        .sel(clk_div),
        .clko(clk_mux2_div)
    );

    wire clk_mux3;
    clkmux_2x1 CLKMUX3 (
        .rst_n(rst_n),
        .clk0(clk_8mhz), 
        .clk1(clk_mux2_div), 
        .sel(sel_mux3),
	    .clko(clk_mux3)
    );

    wire clk_mux4;
    clkmux_2x1 CLKMUX4 (
        .rst_n(rst_n),
        .clk0(clk_8mhz), 
        .clk1(clk_mux3), 
        .sel(sel_mux4),
	    .clko(clk_mux4)
    );

    // Output Clock Divider
    reg     oclkdiv = 0;
    always@(posedge clk_mux4)
        oclkdiv <= oclkdiv + 1'b1;

    wire    clk_mux4_div = oclkdiv;

`ifdef PnR
    (* keep *) sky130_fd_sc_hd__clkbuf_8 clkbuf (
`ifdef USE_POWER_PINS
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPWR),
        .VNB(VGND),
`endif
        .A(clk_mux4),
        .X(clk)
    );
    (* keep *) sky130_fd_sc_hd__clkbuf_8 clk2_buf (
`ifdef USE_POWER_PINS
        .VPWR(VPWR),
        .VGND(VGND),
        .VPB(VPWR),
        .VNB(VGND),
`endif
        .A(clk_mux4_div),
        .X(clk_div_2)
    );
`else // ! PnR
    assign clk = clk_mux4;
    assign clk_div_2 = clk_mux4_div;
`endif // PnR

endmodule
