VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MS_CLK_RST
  CLASS BLOCK ;
  FOREIGN MS_CLK_RST ;
  ORIGIN 0.000 0.000 ;
  SIZE 109.590 BY 120.310 ;
  PIN clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 105.590 78.240 109.590 78.840 ;
    END
  END clk
  PIN clk_div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.747000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END clk_div[0]
  PIN clk_div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.373500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END clk_div[1]
  PIN one
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 116.310 67.990 120.310 ;
    END
  END one
  PIN por_fb_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.576000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 116.310 42.230 120.310 ;
    END
  END por_fb_in
  PIN por_fb_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END por_fb_out
  PIN por_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 105.590 105.440 109.590 106.040 ;
    END
  END por_n
  PIN rst_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END rst_n
  PIN sel_mux0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END sel_mux0
  PIN sel_mux1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 105.590 23.840 109.590 24.440 ;
    END
  END sel_mux1
  PIN sel_mux2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END sel_mux2
  PIN sel_rosc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END sel_rosc[0]
  PIN sel_rosc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 116.310 93.750 120.310 ;
    END
  END sel_rosc[1]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.040 10.640 52.640 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 81.040 10.640 82.640 109.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 36.040 10.640 37.640 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.040 10.640 67.640 109.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 109.040 ;
    END
  END vssd1
  PIN xclk0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END xclk0
  PIN xclk1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END xclk1
  PIN xrst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 116.310 16.470 120.310 ;
    END
  END xrst_n
  PIN zero
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 105.590 51.040 109.590 51.640 ;
    END
  END zero
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 103.960 108.885 ;
      LAYER met1 ;
        RECT 0.070 10.640 104.350 109.040 ;
      LAYER met2 ;
        RECT 0.100 116.030 15.910 116.310 ;
        RECT 16.750 116.030 41.670 116.310 ;
        RECT 42.510 116.030 67.430 116.310 ;
        RECT 68.270 116.030 93.190 116.310 ;
        RECT 94.030 116.030 104.330 116.310 ;
        RECT 0.100 4.280 104.330 116.030 ;
        RECT 0.650 4.000 25.570 4.280 ;
        RECT 26.410 4.000 51.330 4.280 ;
        RECT 52.170 4.000 77.090 4.280 ;
        RECT 77.930 4.000 102.850 4.280 ;
        RECT 103.690 4.000 104.330 4.280 ;
      LAYER met3 ;
        RECT 4.400 108.440 105.590 109.305 ;
        RECT 4.000 106.440 105.590 108.440 ;
        RECT 4.000 105.040 105.190 106.440 ;
        RECT 4.000 82.640 105.590 105.040 ;
        RECT 4.400 81.240 105.590 82.640 ;
        RECT 4.000 79.240 105.590 81.240 ;
        RECT 4.000 77.840 105.190 79.240 ;
        RECT 4.000 55.440 105.590 77.840 ;
        RECT 4.400 54.040 105.590 55.440 ;
        RECT 4.000 52.040 105.590 54.040 ;
        RECT 4.000 50.640 105.190 52.040 ;
        RECT 4.000 28.240 105.590 50.640 ;
        RECT 4.400 26.840 105.590 28.240 ;
        RECT 4.000 24.840 105.590 26.840 ;
        RECT 4.000 23.440 105.190 24.840 ;
        RECT 4.000 10.715 105.590 23.440 ;
  END
END MS_CLK_RST
END LIBRARY

