magic
tech sky130A
magscale 1 2
timestamp 1693328251
<< viali >>
rect 3341 21505 3375 21539
rect 14105 21505 14139 21539
rect 17785 21505 17819 21539
rect 18061 21505 18095 21539
rect 18981 21505 19015 21539
rect 20269 21505 20303 21539
rect 14381 21437 14415 21471
rect 17969 21437 18003 21471
rect 3525 21301 3559 21335
rect 12357 21301 12391 21335
rect 13829 21301 13863 21335
rect 18061 21301 18095 21335
rect 18245 21301 18279 21335
rect 18521 21301 18555 21335
rect 18797 21301 18831 21335
rect 20361 21301 20395 21335
rect 18705 21097 18739 21131
rect 5089 20893 5123 20927
rect 6929 20893 6963 20927
rect 7113 20893 7147 20927
rect 7297 20893 7331 20927
rect 7389 20893 7423 20927
rect 8953 20893 8987 20927
rect 12173 20893 12207 20927
rect 13665 20893 13699 20927
rect 13921 20893 13955 20927
rect 15577 20893 15611 20927
rect 17141 20893 17175 20927
rect 17325 20893 17359 20927
rect 9198 20825 9232 20859
rect 11906 20825 11940 20859
rect 15310 20825 15344 20859
rect 17592 20825 17626 20859
rect 4905 20757 4939 20791
rect 7573 20757 7607 20791
rect 8677 20757 8711 20791
rect 10333 20757 10367 20791
rect 10793 20757 10827 20791
rect 12541 20757 12575 20791
rect 14197 20757 14231 20791
rect 8493 20553 8527 20587
rect 11621 20553 11655 20587
rect 6101 20485 6135 20519
rect 7582 20485 7616 20519
rect 12756 20485 12790 20519
rect 16948 20485 16982 20519
rect 18490 20485 18524 20519
rect 4905 20417 4939 20451
rect 6009 20417 6043 20451
rect 6193 20417 6227 20451
rect 8125 20417 8159 20451
rect 8769 20417 8803 20451
rect 10517 20417 10551 20451
rect 11253 20417 11287 20451
rect 13349 20417 13383 20451
rect 14657 20417 14691 20451
rect 14749 20417 14783 20451
rect 18245 20417 18279 20451
rect 7849 20349 7883 20383
rect 8033 20349 8067 20383
rect 13001 20349 13035 20383
rect 13093 20349 13127 20383
rect 16681 20349 16715 20383
rect 14473 20281 14507 20315
rect 4261 20213 4295 20247
rect 5825 20213 5859 20247
rect 6469 20213 6503 20247
rect 14841 20213 14875 20247
rect 15025 20213 15059 20247
rect 16405 20213 16439 20247
rect 18061 20213 18095 20247
rect 19625 20213 19659 20247
rect 7297 20009 7331 20043
rect 10333 20009 10367 20043
rect 12909 20009 12943 20043
rect 14289 20009 14323 20043
rect 16957 20009 16991 20043
rect 17417 20009 17451 20043
rect 17693 20009 17727 20043
rect 10517 19873 10551 19907
rect 19073 19873 19107 19907
rect 4077 19805 4111 19839
rect 6285 19805 6319 19839
rect 6469 19805 6503 19839
rect 7113 19805 7147 19839
rect 10784 19805 10818 19839
rect 15577 19805 15611 19839
rect 18806 19805 18840 19839
rect 6929 19737 6963 19771
rect 12081 19737 12115 19771
rect 12357 19737 12391 19771
rect 12633 19737 12667 19771
rect 14473 19737 14507 19771
rect 15844 19737 15878 19771
rect 4077 19669 4111 19703
rect 6377 19669 6411 19703
rect 11897 19669 11931 19703
rect 12265 19669 12299 19703
rect 12449 19669 12483 19703
rect 14105 19669 14139 19703
rect 14268 19669 14302 19703
rect 15393 19669 15427 19703
rect 6094 19465 6128 19499
rect 10057 19465 10091 19499
rect 11345 19465 11379 19499
rect 15025 19465 15059 19499
rect 17877 19465 17911 19499
rect 17969 19465 18003 19499
rect 18061 19465 18095 19499
rect 7582 19397 7616 19431
rect 12734 19397 12768 19431
rect 14197 19397 14231 19431
rect 14413 19397 14447 19431
rect 18245 19397 18279 19431
rect 18889 19397 18923 19431
rect 20186 19397 20220 19431
rect 2513 19329 2547 19363
rect 3157 19329 3191 19363
rect 3249 19329 3283 19363
rect 4620 19329 4654 19363
rect 5917 19329 5951 19363
rect 6009 19329 6043 19363
rect 6193 19329 6227 19363
rect 8309 19329 8343 19363
rect 10885 19329 10919 19363
rect 11069 19329 11103 19363
rect 11161 19329 11195 19363
rect 13001 19329 13035 19363
rect 14657 19329 14691 19363
rect 14841 19329 14875 19363
rect 20453 19329 20487 19363
rect 4353 19261 4387 19295
rect 7849 19261 7883 19295
rect 8125 19261 8159 19295
rect 8585 19261 8619 19295
rect 6469 19193 6503 19227
rect 14565 19193 14599 19227
rect 3249 19125 3283 19159
rect 4169 19125 4203 19159
rect 5733 19125 5767 19159
rect 10793 19125 10827 19159
rect 11161 19125 11195 19159
rect 11621 19125 11655 19159
rect 14381 19125 14415 19159
rect 14657 19125 14691 19159
rect 17693 19125 17727 19159
rect 19073 19125 19107 19159
rect 4537 18921 4571 18955
rect 6285 18921 6319 18955
rect 6469 18921 6503 18955
rect 9045 18921 9079 18955
rect 11253 18921 11287 18955
rect 13829 18921 13863 18955
rect 15301 18921 15335 18955
rect 16957 18921 16991 18955
rect 18337 18921 18371 18955
rect 19625 18921 19659 18955
rect 6745 18853 6779 18887
rect 7849 18853 7883 18887
rect 12817 18853 12851 18887
rect 17325 18853 17359 18887
rect 4997 18785 5031 18819
rect 11437 18785 11471 18819
rect 14657 18785 14691 18819
rect 15393 18785 15427 18819
rect 17049 18785 17083 18819
rect 18429 18785 18463 18819
rect 19625 18785 19659 18819
rect 1961 18717 1995 18751
rect 2605 18717 2639 18751
rect 2697 18717 2731 18751
rect 4905 18717 4939 18751
rect 9137 18717 9171 18751
rect 15649 18717 15683 18751
rect 16957 18717 16991 18751
rect 18521 18717 18555 18751
rect 19441 18717 19475 18751
rect 19717 18717 19751 18751
rect 6101 18649 6135 18683
rect 11704 18649 11738 18683
rect 14105 18649 14139 18683
rect 2881 18581 2915 18615
rect 6301 18581 6335 18615
rect 14289 18581 14323 18615
rect 14381 18581 14415 18615
rect 14473 18581 14507 18615
rect 16773 18581 16807 18615
rect 18153 18581 18187 18615
rect 19257 18581 19291 18615
rect 12265 18377 12299 18411
rect 13737 18377 13771 18411
rect 15945 18377 15979 18411
rect 16773 18377 16807 18411
rect 19625 18377 19659 18411
rect 12624 18309 12658 18343
rect 15485 18309 15519 18343
rect 16129 18309 16163 18343
rect 16345 18309 16379 18343
rect 17886 18309 17920 18343
rect 18512 18309 18546 18343
rect 7573 18241 7607 18275
rect 8033 18241 8067 18275
rect 12357 18241 12391 18275
rect 15126 18241 15160 18275
rect 15761 18241 15795 18275
rect 18153 18241 18187 18275
rect 18245 18241 18279 18275
rect 4721 18173 4755 18207
rect 7665 18173 7699 18207
rect 8309 18173 8343 18207
rect 15393 18173 15427 18207
rect 15577 18173 15611 18207
rect 7941 18105 7975 18139
rect 9781 18037 9815 18071
rect 14013 18037 14047 18071
rect 15577 18037 15611 18071
rect 16313 18037 16347 18071
rect 16497 18037 16531 18071
rect 9689 17833 9723 17867
rect 13829 17833 13863 17867
rect 14197 17833 14231 17867
rect 15853 17833 15887 17867
rect 18061 17833 18095 17867
rect 9413 17765 9447 17799
rect 1685 17697 1719 17731
rect 1961 17697 1995 17731
rect 4169 17697 4203 17731
rect 5641 17697 5675 17731
rect 6101 17697 6135 17731
rect 15577 17697 15611 17731
rect 18521 17697 18555 17731
rect 1593 17629 1627 17663
rect 3893 17629 3927 17663
rect 5825 17629 5859 17663
rect 8585 17629 8619 17663
rect 8769 17629 8803 17663
rect 9137 17629 9171 17663
rect 9413 17629 9447 17663
rect 10333 17629 10367 17663
rect 15310 17629 15344 17663
rect 16966 17629 17000 17663
rect 17233 17629 17267 17663
rect 19533 17629 19567 17663
rect 19625 17629 19659 17663
rect 9673 17561 9707 17595
rect 9873 17561 9907 17595
rect 9965 17561 9999 17595
rect 10149 17561 10183 17595
rect 10241 17561 10275 17595
rect 17877 17561 17911 17595
rect 18093 17561 18127 17595
rect 19257 17561 19291 17595
rect 19441 17561 19475 17595
rect 19809 17561 19843 17595
rect 2973 17493 3007 17527
rect 3249 17493 3283 17527
rect 7573 17493 7607 17527
rect 8677 17493 8711 17527
rect 9229 17493 9263 17527
rect 9505 17493 9539 17527
rect 10517 17493 10551 17527
rect 18245 17493 18279 17527
rect 5181 17289 5215 17323
rect 10517 17289 10551 17323
rect 12541 17289 12575 17323
rect 15577 17289 15611 17323
rect 16865 17289 16899 17323
rect 18061 17289 18095 17323
rect 3516 17221 3550 17255
rect 9045 17221 9079 17255
rect 10977 17221 11011 17255
rect 13952 17221 13986 17255
rect 19472 17221 19506 17255
rect 1685 17153 1719 17187
rect 1952 17153 1986 17187
rect 4997 17153 5031 17187
rect 5365 17153 5399 17187
rect 5549 17153 5583 17187
rect 5641 17153 5675 17187
rect 5825 17153 5859 17187
rect 10609 17153 10643 17187
rect 10793 17153 10827 17187
rect 10885 17153 10919 17187
rect 11069 17153 11103 17187
rect 14197 17153 14231 17187
rect 19717 17153 19751 17187
rect 3249 17085 3283 17119
rect 4813 17085 4847 17119
rect 5733 17085 5767 17119
rect 6837 17085 6871 17119
rect 7113 17085 7147 17119
rect 8769 17085 8803 17119
rect 3065 16949 3099 16983
rect 4629 16949 4663 16983
rect 5549 16949 5583 16983
rect 8585 16949 8619 16983
rect 10793 16949 10827 16983
rect 12817 16949 12851 16983
rect 18337 16949 18371 16983
rect 3985 16745 4019 16779
rect 4169 16745 4203 16779
rect 5641 16745 5675 16779
rect 10866 16745 10900 16779
rect 12357 16745 12391 16779
rect 14381 16745 14415 16779
rect 17417 16745 17451 16779
rect 3433 16677 3467 16711
rect 4537 16677 4571 16711
rect 1685 16609 1719 16643
rect 1869 16609 1903 16643
rect 5733 16609 5767 16643
rect 8677 16609 8711 16643
rect 10517 16609 10551 16643
rect 10609 16609 10643 16643
rect 15117 16609 15151 16643
rect 15393 16609 15427 16643
rect 15577 16609 15611 16643
rect 15853 16609 15887 16643
rect 17601 16609 17635 16643
rect 2136 16541 2170 16575
rect 3433 16541 3467 16575
rect 3617 16541 3651 16575
rect 4261 16541 4295 16575
rect 5989 16541 6023 16575
rect 14565 16541 14599 16575
rect 15209 16541 15243 16575
rect 15669 16541 15703 16575
rect 17868 16541 17902 16575
rect 1501 16473 1535 16507
rect 3801 16473 3835 16507
rect 4353 16473 4387 16507
rect 4537 16473 4571 16507
rect 14933 16473 14967 16507
rect 15301 16473 15335 16507
rect 3249 16405 3283 16439
rect 4001 16405 4035 16439
rect 7113 16405 7147 16439
rect 14749 16405 14783 16439
rect 14841 16405 14875 16439
rect 18981 16405 19015 16439
rect 1961 16201 1995 16235
rect 12725 16201 12759 16235
rect 14289 16201 14323 16235
rect 16405 16201 16439 16235
rect 13154 16133 13188 16167
rect 14473 16133 14507 16167
rect 17233 16133 17267 16167
rect 17601 16133 17635 16167
rect 18429 16133 18463 16167
rect 2053 16065 2087 16099
rect 10333 16065 10367 16099
rect 10517 16065 10551 16099
rect 12909 16065 12943 16099
rect 14657 16065 14691 16099
rect 14749 16065 14783 16099
rect 15281 16065 15315 16099
rect 17969 16065 18003 16099
rect 18061 16065 18095 16099
rect 20094 16065 20128 16099
rect 20361 16065 20395 16099
rect 15025 15997 15059 16031
rect 18245 15997 18279 16031
rect 18337 15997 18371 16031
rect 17325 15929 17359 15963
rect 17601 15929 17635 15963
rect 3525 15861 3559 15895
rect 10425 15861 10459 15895
rect 11069 15861 11103 15895
rect 14657 15861 14691 15895
rect 14933 15861 14967 15895
rect 17417 15861 17451 15895
rect 17785 15861 17819 15895
rect 18705 15861 18739 15895
rect 18981 15861 19015 15895
rect 13829 15657 13863 15691
rect 15853 15657 15887 15691
rect 15945 15657 15979 15691
rect 16957 15657 16991 15691
rect 18613 15657 18647 15691
rect 18889 15657 18923 15691
rect 20453 15657 20487 15691
rect 4353 15589 4387 15623
rect 15485 15589 15519 15623
rect 15669 15589 15703 15623
rect 19809 15589 19843 15623
rect 6377 15521 6411 15555
rect 9965 15521 9999 15555
rect 10517 15521 10551 15555
rect 14105 15521 14139 15555
rect 16037 15521 16071 15555
rect 19257 15521 19291 15555
rect 3801 15453 3835 15487
rect 4077 15453 4111 15487
rect 4169 15453 4203 15487
rect 4445 15453 4479 15487
rect 4905 15453 4939 15487
rect 9413 15453 9447 15487
rect 9505 15453 9539 15487
rect 9689 15453 9723 15487
rect 9873 15453 9907 15487
rect 10609 15453 10643 15487
rect 11161 15453 11195 15487
rect 14372 15453 14406 15487
rect 15669 15453 15703 15487
rect 18337 15453 18371 15487
rect 18797 15453 18831 15487
rect 18889 15453 18923 15487
rect 19073 15453 19107 15487
rect 19625 15453 19659 15487
rect 20269 15453 20303 15487
rect 3985 15385 4019 15419
rect 4537 15385 4571 15419
rect 6653 15385 6687 15419
rect 10149 15385 10183 15419
rect 10333 15385 10367 15419
rect 11437 15385 11471 15419
rect 13001 15385 13035 15419
rect 13369 15385 13403 15419
rect 18092 15385 18126 15419
rect 4721 15317 4755 15351
rect 8125 15317 8159 15351
rect 9229 15317 9263 15351
rect 10977 15317 11011 15351
rect 12909 15317 12943 15351
rect 16681 15317 16715 15351
rect 19441 15317 19475 15351
rect 19533 15317 19567 15351
rect 3801 15113 3835 15147
rect 4353 15113 4387 15147
rect 6653 15113 6687 15147
rect 12081 15113 12115 15147
rect 14105 15113 14139 15147
rect 14381 15113 14415 15147
rect 17141 15113 17175 15147
rect 17325 15113 17359 15147
rect 18521 15113 18555 15147
rect 1869 15045 1903 15079
rect 2329 15045 2363 15079
rect 3893 15045 3927 15079
rect 7021 15045 7055 15079
rect 8861 15045 8895 15079
rect 11805 15045 11839 15079
rect 15494 15045 15528 15079
rect 18245 15045 18279 15079
rect 1501 14977 1535 15011
rect 1685 14977 1719 15011
rect 1777 14977 1811 15011
rect 6469 14977 6503 15011
rect 8585 14977 8619 15011
rect 10885 14977 10919 15011
rect 11069 14977 11103 15011
rect 11713 14977 11747 15011
rect 11897 14977 11931 15011
rect 12633 14977 12667 15011
rect 15761 14977 15795 15011
rect 17233 14977 17267 15011
rect 17509 14977 17543 15011
rect 17601 14977 17635 15011
rect 19634 14977 19668 15011
rect 19901 14977 19935 15011
rect 2053 14909 2087 14943
rect 4445 14909 4479 14943
rect 5917 14909 5951 14943
rect 6193 14909 6227 14943
rect 6745 14909 6779 14943
rect 10333 14909 10367 14943
rect 10977 14909 11011 14943
rect 11160 14909 11194 14943
rect 11345 14909 11379 14943
rect 4169 14841 4203 14875
rect 11529 14841 11563 14875
rect 12265 14841 12299 14875
rect 16957 14841 16991 14875
rect 17785 14841 17819 14875
rect 1501 14773 1535 14807
rect 8493 14773 8527 14807
rect 12173 14773 12207 14807
rect 3157 14569 3191 14603
rect 5549 14569 5583 14603
rect 6745 14569 6779 14603
rect 7481 14569 7515 14603
rect 8493 14569 8527 14603
rect 6929 14501 6963 14535
rect 7113 14501 7147 14535
rect 14749 14501 14783 14535
rect 1685 14433 1719 14467
rect 3801 14433 3835 14467
rect 4077 14433 4111 14467
rect 13185 14433 13219 14467
rect 14933 14433 14967 14467
rect 1409 14365 1443 14399
rect 6653 14365 6687 14399
rect 7481 14365 7515 14399
rect 7665 14365 7699 14399
rect 11161 14365 11195 14399
rect 11437 14365 11471 14399
rect 7389 14297 7423 14331
rect 11713 14297 11747 14331
rect 15200 14297 15234 14331
rect 11069 14229 11103 14263
rect 11345 14229 11379 14263
rect 16313 14229 16347 14263
rect 16681 14229 16715 14263
rect 9137 14025 9171 14059
rect 14105 14025 14139 14059
rect 14381 14025 14415 14059
rect 16313 14025 16347 14059
rect 18521 14025 18555 14059
rect 18797 14025 18831 14059
rect 7113 13957 7147 13991
rect 15516 13957 15550 13991
rect 15853 13957 15887 13991
rect 19910 13957 19944 13991
rect 2237 13889 2271 13923
rect 6924 13889 6958 13923
rect 7021 13889 7055 13923
rect 7297 13889 7331 13923
rect 8677 13889 8711 13923
rect 8953 13889 8987 13923
rect 10057 13889 10091 13923
rect 16129 13889 16163 13923
rect 16937 13889 16971 13923
rect 20177 13889 20211 13923
rect 2145 13821 2179 13855
rect 10517 13821 10551 13855
rect 11069 13821 11103 13855
rect 15761 13821 15795 13855
rect 15945 13821 15979 13855
rect 16681 13821 16715 13855
rect 6745 13685 6779 13719
rect 8769 13685 8803 13719
rect 10149 13685 10183 13719
rect 15945 13685 15979 13719
rect 18061 13685 18095 13719
rect 5076 13481 5110 13515
rect 8401 13481 8435 13515
rect 11345 13481 11379 13515
rect 3157 13413 3191 13447
rect 4629 13413 4663 13447
rect 15485 13413 15519 13447
rect 17049 13413 17083 13447
rect 1409 13345 1443 13379
rect 4813 13345 4847 13379
rect 8953 13345 8987 13379
rect 13185 13345 13219 13379
rect 13829 13345 13863 13379
rect 14105 13345 14139 13379
rect 4077 13277 4111 13311
rect 4353 13277 4387 13311
rect 4497 13277 4531 13311
rect 6653 13277 6687 13311
rect 10793 13277 10827 13311
rect 11213 13277 11247 13311
rect 15669 13277 15703 13311
rect 15936 13277 15970 13311
rect 17417 13277 17451 13311
rect 19073 13277 19107 13311
rect 1685 13209 1719 13243
rect 3525 13209 3559 13243
rect 4261 13209 4295 13243
rect 6929 13209 6963 13243
rect 8677 13209 8711 13243
rect 9229 13209 9263 13243
rect 10977 13209 11011 13243
rect 11069 13209 11103 13243
rect 14372 13209 14406 13243
rect 18806 13209 18840 13243
rect 6561 13141 6595 13175
rect 8585 13141 8619 13175
rect 10701 13141 10735 13175
rect 17693 13141 17727 13175
rect 2237 12937 2271 12971
rect 4353 12937 4387 12971
rect 6193 12937 6227 12971
rect 6561 12937 6595 12971
rect 9505 12937 9539 12971
rect 11345 12937 11379 12971
rect 13277 12937 13311 12971
rect 14749 12937 14783 12971
rect 15761 12937 15795 12971
rect 15853 12937 15887 12971
rect 15945 12937 15979 12971
rect 17601 12937 17635 12971
rect 19349 12937 19383 12971
rect 4721 12869 4755 12903
rect 11805 12869 11839 12903
rect 16129 12869 16163 12903
rect 17325 12869 17359 12903
rect 1685 12801 1719 12835
rect 2421 12801 2455 12835
rect 6469 12801 6503 12835
rect 7757 12801 7791 12835
rect 9597 12801 9631 12835
rect 13369 12801 13403 12835
rect 13636 12801 13670 12835
rect 15485 12801 15519 12835
rect 17509 12801 17543 12835
rect 17693 12801 17727 12835
rect 18236 12801 18270 12835
rect 2145 12733 2179 12767
rect 2605 12733 2639 12767
rect 2881 12733 2915 12767
rect 4445 12733 4479 12767
rect 8033 12733 8067 12767
rect 9873 12733 9907 12767
rect 11529 12733 11563 12767
rect 17969 12733 18003 12767
rect 2053 12665 2087 12699
rect 15577 12597 15611 12631
rect 17141 12597 17175 12631
rect 17877 12597 17911 12631
rect 3801 12393 3835 12427
rect 4721 12393 4755 12427
rect 8493 12393 8527 12427
rect 9965 12393 9999 12427
rect 11161 12393 11195 12427
rect 12357 12393 12391 12427
rect 13829 12393 13863 12427
rect 14657 12393 14691 12427
rect 16037 12393 16071 12427
rect 16313 12393 16347 12427
rect 18889 12393 18923 12427
rect 10977 12325 11011 12359
rect 14105 12325 14139 12359
rect 2145 12257 2179 12291
rect 3617 12257 3651 12291
rect 16957 12257 16991 12291
rect 18889 12257 18923 12291
rect 1869 12189 1903 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 4537 12189 4571 12223
rect 4813 12189 4847 12223
rect 8309 12189 8343 12223
rect 8493 12189 8527 12223
rect 8953 12189 8987 12223
rect 9045 12189 9079 12223
rect 9781 12189 9815 12223
rect 9965 12189 9999 12223
rect 10885 12189 10919 12223
rect 11345 12189 11379 12223
rect 12449 12189 12483 12223
rect 14289 12189 14323 12223
rect 16313 12189 16347 12223
rect 16405 12189 16439 12223
rect 17224 12189 17258 12223
rect 18705 12189 18739 12223
rect 18981 12189 19015 12223
rect 12694 12121 12728 12155
rect 15853 12121 15887 12155
rect 16053 12121 16087 12155
rect 14381 12053 14415 12087
rect 14473 12053 14507 12087
rect 16221 12053 16255 12087
rect 16681 12053 16715 12087
rect 18337 12053 18371 12087
rect 18521 12053 18555 12087
rect 1593 11849 1627 11883
rect 2513 11849 2547 11883
rect 4353 11849 4387 11883
rect 14289 11849 14323 11883
rect 15685 11849 15719 11883
rect 15853 11849 15887 11883
rect 16313 11849 16347 11883
rect 18153 11849 18187 11883
rect 18889 11849 18923 11883
rect 13829 11781 13863 11815
rect 15485 11781 15519 11815
rect 16957 11781 16991 11815
rect 17325 11781 17359 11815
rect 18061 11781 18095 11815
rect 20002 11781 20036 11815
rect 1409 11713 1443 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 15945 11713 15979 11747
rect 17509 11713 17543 11747
rect 18337 11713 18371 11747
rect 20269 11713 20303 11747
rect 16037 11645 16071 11679
rect 17601 11645 17635 11679
rect 17785 11645 17819 11679
rect 17877 11645 17911 11679
rect 17969 11645 18003 11679
rect 18245 11645 18279 11679
rect 18429 11645 18463 11679
rect 13921 11509 13955 11543
rect 15669 11509 15703 11543
rect 16129 11509 16163 11543
rect 9137 11305 9171 11339
rect 9597 11305 9631 11339
rect 11897 11305 11931 11339
rect 12357 11305 12391 11339
rect 12541 11305 12575 11339
rect 9321 11237 9355 11271
rect 9689 11237 9723 11271
rect 4445 11169 4479 11203
rect 10241 11169 10275 11203
rect 10885 11169 10919 11203
rect 11345 11169 11379 11203
rect 16681 11169 16715 11203
rect 18613 11169 18647 11203
rect 18981 11169 19015 11203
rect 1593 11101 1627 11135
rect 2237 11101 2271 11135
rect 2329 11101 2363 11135
rect 2881 11101 2915 11135
rect 6285 11101 6319 11135
rect 8493 11101 8527 11135
rect 9413 11101 9447 11135
rect 10425 11101 10459 11135
rect 10701 11101 10735 11135
rect 10977 11101 11011 11135
rect 11437 11101 11471 11135
rect 13665 11101 13699 11135
rect 13921 11101 13955 11135
rect 3985 11033 4019 11067
rect 4169 11033 4203 11067
rect 4721 11033 4755 11067
rect 6653 11033 6687 11067
rect 8953 11033 8987 11067
rect 9153 11033 9187 11067
rect 9873 11033 9907 11067
rect 10057 11033 10091 11067
rect 10609 11033 10643 11067
rect 16414 11033 16448 11067
rect 2513 10965 2547 10999
rect 2697 10965 2731 10999
rect 4353 10965 4387 10999
rect 6193 10965 6227 10999
rect 8309 10965 8343 10999
rect 11621 10965 11655 10999
rect 14749 10965 14783 10999
rect 15025 10965 15059 10999
rect 15301 10965 15335 10999
rect 4077 10761 4111 10795
rect 5181 10761 5215 10795
rect 9459 10761 9493 10795
rect 9873 10761 9907 10795
rect 10057 10761 10091 10795
rect 11161 10761 11195 10795
rect 13461 10761 13495 10795
rect 16313 10761 16347 10795
rect 16957 10761 16991 10795
rect 18429 10761 18463 10795
rect 4997 10693 5031 10727
rect 5733 10693 5767 10727
rect 11805 10693 11839 10727
rect 14596 10693 14630 10727
rect 19818 10693 19852 10727
rect 2237 10625 2271 10659
rect 2329 10625 2363 10659
rect 4353 10625 4387 10659
rect 4445 10625 4479 10659
rect 4537 10625 4571 10659
rect 4655 10625 4689 10659
rect 4905 10625 4939 10659
rect 5089 10625 5123 10659
rect 5365 10625 5399 10659
rect 5457 10625 5491 10659
rect 6193 10625 6227 10659
rect 6377 10625 6411 10659
rect 6561 10625 6595 10659
rect 6653 10625 6687 10659
rect 6745 10625 6779 10659
rect 7573 10625 7607 10659
rect 11529 10625 11563 10659
rect 14841 10625 14875 10659
rect 14933 10625 14967 10659
rect 15200 10625 15234 10659
rect 17049 10625 17083 10659
rect 17316 10625 17350 10659
rect 20085 10625 20119 10659
rect 2605 10557 2639 10591
rect 4169 10557 4203 10591
rect 4813 10557 4847 10591
rect 5825 10557 5859 10591
rect 5917 10557 5951 10591
rect 7665 10557 7699 10591
rect 8033 10557 8067 10591
rect 10517 10557 10551 10591
rect 13277 10557 13311 10591
rect 6009 10489 6043 10523
rect 10425 10489 10459 10523
rect 1593 10421 1627 10455
rect 6101 10421 6135 10455
rect 6929 10421 6963 10455
rect 10057 10421 10091 10455
rect 18705 10421 18739 10455
rect 2132 10217 2166 10251
rect 3801 10217 3835 10251
rect 4905 10217 4939 10251
rect 5089 10217 5123 10251
rect 5549 10217 5583 10251
rect 5917 10217 5951 10251
rect 6101 10217 6135 10251
rect 8401 10217 8435 10251
rect 9505 10217 9539 10251
rect 15485 10217 15519 10251
rect 16497 10217 16531 10251
rect 18245 10217 18279 10251
rect 6285 10149 6319 10183
rect 9321 10149 9355 10183
rect 1869 10081 1903 10115
rect 4353 10081 4387 10115
rect 5733 10081 5767 10115
rect 7757 10081 7791 10115
rect 10057 10081 10091 10115
rect 11897 10081 11931 10115
rect 13277 10081 13311 10115
rect 13921 10081 13955 10115
rect 14105 10081 14139 10115
rect 16589 10081 16623 10115
rect 18521 10081 18555 10115
rect 18705 10081 18739 10115
rect 20453 10081 20487 10115
rect 1593 10013 1627 10047
rect 4261 10013 4295 10047
rect 5641 10013 5675 10047
rect 5917 10013 5951 10047
rect 8033 10013 8067 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 9689 10013 9723 10047
rect 16856 10013 16890 10047
rect 18429 10013 18463 10047
rect 20177 10013 20211 10047
rect 4721 9945 4755 9979
rect 4937 9945 4971 9979
rect 5181 9945 5215 9979
rect 5365 9945 5399 9979
rect 8585 9945 8619 9979
rect 8769 9945 8803 9979
rect 8953 9945 8987 9979
rect 11621 9945 11655 9979
rect 14372 9945 14406 9979
rect 18797 9945 18831 9979
rect 18889 9945 18923 9979
rect 1685 9877 1719 9911
rect 3617 9877 3651 9911
rect 4169 9877 4203 9911
rect 10149 9877 10183 9911
rect 17969 9877 18003 9911
rect 2513 9673 2547 9707
rect 6469 9673 6503 9707
rect 7757 9673 7791 9707
rect 8125 9673 8159 9707
rect 10333 9673 10367 9707
rect 15485 9673 15519 9707
rect 17509 9673 17543 9707
rect 3801 9605 3835 9639
rect 6193 9605 6227 9639
rect 17785 9605 17819 9639
rect 1593 9537 1627 9571
rect 6377 9537 6411 9571
rect 6561 9537 6595 9571
rect 6745 9537 6779 9571
rect 6929 9537 6963 9571
rect 7941 9537 7975 9571
rect 8033 9537 8067 9571
rect 8401 9537 8435 9571
rect 8585 9537 8619 9571
rect 17417 9537 17451 9571
rect 17693 9537 17727 9571
rect 18153 9537 18187 9571
rect 18429 9537 18463 9571
rect 19726 9537 19760 9571
rect 19993 9537 20027 9571
rect 8263 9469 8297 9503
rect 8861 9469 8895 9503
rect 18245 9469 18279 9503
rect 17601 9401 17635 9435
rect 17969 9401 18003 9435
rect 18613 9401 18647 9435
rect 2237 9333 2271 9367
rect 6745 9333 6779 9367
rect 8401 9333 8435 9367
rect 18429 9333 18463 9367
rect 6285 9129 6319 9163
rect 8769 9129 8803 9163
rect 17417 9129 17451 9163
rect 17785 9129 17819 9163
rect 19073 9129 19107 9163
rect 18337 9061 18371 9095
rect 17141 8993 17175 9027
rect 2329 8925 2363 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 7113 8925 7147 8959
rect 7389 8925 7423 8959
rect 7849 8925 7883 8959
rect 8493 8925 8527 8959
rect 8769 8925 8803 8959
rect 10609 8925 10643 8959
rect 13921 8925 13955 8959
rect 14105 8925 14139 8959
rect 14372 8925 14406 8959
rect 17601 8925 17635 8959
rect 17785 8925 17819 8959
rect 18705 8925 18739 8959
rect 4905 8857 4939 8891
rect 10885 8857 10919 8891
rect 16874 8857 16908 8891
rect 18521 8857 18555 8891
rect 1685 8789 1719 8823
rect 4537 8789 4571 8823
rect 6929 8789 6963 8823
rect 7297 8789 7331 8823
rect 7757 8789 7791 8823
rect 8585 8789 8619 8823
rect 12357 8789 12391 8823
rect 15485 8789 15519 8823
rect 15761 8789 15795 8823
rect 18797 8789 18831 8823
rect 18889 8789 18923 8823
rect 3709 8585 3743 8619
rect 5365 8585 5399 8619
rect 5641 8585 5675 8619
rect 10517 8585 10551 8619
rect 11261 8585 11295 8619
rect 16329 8585 16363 8619
rect 16497 8585 16531 8619
rect 17049 8585 17083 8619
rect 4169 8517 4203 8551
rect 4261 8517 4295 8551
rect 4997 8517 5031 8551
rect 9321 8517 9355 8551
rect 10885 8517 10919 8551
rect 16129 8517 16163 8551
rect 17233 8517 17267 8551
rect 17449 8517 17483 8551
rect 1685 8449 1719 8483
rect 4077 8449 4111 8483
rect 4379 8449 4413 8483
rect 4629 8449 4663 8483
rect 4721 8449 4755 8483
rect 4905 8449 4939 8483
rect 5181 8449 5215 8483
rect 5273 8449 5307 8483
rect 5825 8449 5859 8483
rect 6101 8449 6135 8483
rect 6469 8449 6503 8483
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 10701 8449 10735 8483
rect 10977 8449 11011 8483
rect 11121 8449 11155 8483
rect 11713 8449 11747 8483
rect 16681 8449 16715 8483
rect 17877 8449 17911 8483
rect 18144 8449 18178 8483
rect 4537 8381 4571 8415
rect 5917 8381 5951 8415
rect 6745 8381 6779 8415
rect 8953 8381 8987 8415
rect 11989 8381 12023 8415
rect 13829 8381 13863 8415
rect 15577 8381 15611 8415
rect 16773 8381 16807 8415
rect 8401 8313 8435 8347
rect 9689 8313 9723 8347
rect 17601 8313 17635 8347
rect 19257 8313 19291 8347
rect 2421 8245 2455 8279
rect 3893 8245 3927 8279
rect 4813 8245 4847 8279
rect 5549 8245 5583 8279
rect 5825 8245 5859 8279
rect 8217 8245 8251 8279
rect 9137 8245 9171 8279
rect 9321 8245 9355 8279
rect 11897 8245 11931 8279
rect 12246 8245 12280 8279
rect 13737 8245 13771 8279
rect 14086 8245 14120 8279
rect 16313 8245 16347 8279
rect 16865 8245 16899 8279
rect 17417 8245 17451 8279
rect 2132 8041 2166 8075
rect 5549 8041 5583 8075
rect 7297 8041 7331 8075
rect 7573 8041 7607 8075
rect 7757 8041 7791 8075
rect 8217 8041 8251 8075
rect 11529 8041 11563 8075
rect 13737 8041 13771 8075
rect 16129 8041 16163 8075
rect 17693 8041 17727 8075
rect 19257 8041 19291 8075
rect 20177 8041 20211 8075
rect 20361 8041 20395 8075
rect 11345 7973 11379 8007
rect 17141 7973 17175 8007
rect 17509 7973 17543 8007
rect 19809 7973 19843 8007
rect 1869 7905 1903 7939
rect 3801 7905 3835 7939
rect 6377 7905 6411 7939
rect 6653 7905 6687 7939
rect 8677 7905 8711 7939
rect 8953 7905 8987 7939
rect 10701 7905 10735 7939
rect 12081 7905 12115 7939
rect 19993 7905 20027 7939
rect 5641 7837 5675 7871
rect 5825 7837 5859 7871
rect 6009 7837 6043 7871
rect 6285 7837 6319 7871
rect 6469 7837 6503 7871
rect 7021 7837 7055 7871
rect 7113 7837 7147 7871
rect 11805 7837 11839 7871
rect 13645 7837 13679 7871
rect 14749 7837 14783 7871
rect 15016 7837 15050 7871
rect 19073 7837 19107 7871
rect 19441 7837 19475 7871
rect 19901 7837 19935 7871
rect 20177 7837 20211 7871
rect 4077 7769 4111 7803
rect 5917 7769 5951 7803
rect 6791 7769 6825 7803
rect 6929 7769 6963 7803
rect 7389 7769 7423 7803
rect 8401 7769 8435 7803
rect 10425 7769 10459 7803
rect 11069 7769 11103 7803
rect 18828 7769 18862 7803
rect 3617 7701 3651 7735
rect 6193 7701 6227 7735
rect 7599 7701 7633 7735
rect 13553 7701 13587 7735
rect 14657 7701 14691 7735
rect 19533 7701 19567 7735
rect 19625 7701 19659 7735
rect 3709 7497 3743 7531
rect 4537 7497 4571 7531
rect 5733 7497 5767 7531
rect 8585 7497 8619 7531
rect 11621 7497 11655 7531
rect 18613 7497 18647 7531
rect 2421 7429 2455 7463
rect 4905 7429 4939 7463
rect 5273 7429 5307 7463
rect 6653 7429 6687 7463
rect 10149 7429 10183 7463
rect 15200 7429 15234 7463
rect 18429 7429 18463 7463
rect 4721 7361 4755 7395
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 5181 7361 5215 7395
rect 5365 7361 5399 7395
rect 5457 7361 5491 7395
rect 5641 7361 5675 7395
rect 6377 7361 6411 7395
rect 8769 7361 8803 7395
rect 9229 7361 9263 7395
rect 9321 7361 9355 7395
rect 9505 7361 9539 7395
rect 11529 7361 11563 7395
rect 14841 7361 14875 7395
rect 14933 7361 14967 7395
rect 19726 7361 19760 7395
rect 19993 7361 20027 7395
rect 1593 7293 1627 7327
rect 8861 7293 8895 7327
rect 5917 7157 5951 7191
rect 8125 7157 8159 7191
rect 10057 7157 10091 7191
rect 16313 7157 16347 7191
rect 6285 6953 6319 6987
rect 17509 6953 17543 6987
rect 17693 6953 17727 6987
rect 18429 6953 18463 6987
rect 16957 6885 16991 6919
rect 2237 6817 2271 6851
rect 12817 6749 12851 6783
rect 15301 6749 15335 6783
rect 15393 6749 15427 6783
rect 15660 6749 15694 6783
rect 17785 6749 17819 6783
rect 17877 6749 17911 6783
rect 1501 6681 1535 6715
rect 17233 6681 17267 6715
rect 17325 6681 17359 6715
rect 17601 6681 17635 6715
rect 12909 6613 12943 6647
rect 16773 6613 16807 6647
rect 17141 6613 17175 6647
rect 18061 6613 18095 6647
rect 7573 6409 7607 6443
rect 9505 6409 9539 6443
rect 14105 6409 14139 6443
rect 18061 6409 18095 6443
rect 14473 6341 14507 6375
rect 18490 6341 18524 6375
rect 2789 6273 2823 6307
rect 3065 6273 3099 6307
rect 7757 6273 7791 6307
rect 10977 6273 11011 6307
rect 12357 6273 12391 6307
rect 14197 6273 14231 6307
rect 16937 6273 16971 6307
rect 18245 6273 18279 6307
rect 8033 6205 8067 6239
rect 11069 6205 11103 6239
rect 12633 6205 12667 6239
rect 16497 6205 16531 6239
rect 16681 6205 16715 6239
rect 2605 6069 2639 6103
rect 3157 6069 3191 6103
rect 10701 6069 10735 6103
rect 15945 6069 15979 6103
rect 19625 6069 19659 6103
rect 6101 5865 6135 5899
rect 7941 5865 7975 5899
rect 12449 5865 12483 5899
rect 13093 5865 13127 5899
rect 16589 5865 16623 5899
rect 16773 5865 16807 5899
rect 11437 5797 11471 5831
rect 1869 5729 1903 5763
rect 2145 5729 2179 5763
rect 3617 5729 3651 5763
rect 4077 5729 4111 5763
rect 6193 5729 6227 5763
rect 11897 5729 11931 5763
rect 12081 5729 12115 5763
rect 18153 5729 18187 5763
rect 1409 5661 1443 5695
rect 3801 5661 3835 5695
rect 8033 5661 8067 5695
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 9781 5661 9815 5695
rect 10057 5661 10091 5695
rect 10324 5661 10358 5695
rect 11713 5661 11747 5695
rect 11989 5661 12023 5695
rect 12173 5661 12207 5695
rect 12633 5661 12667 5695
rect 12817 5661 12851 5695
rect 13001 5661 13035 5695
rect 13277 5661 13311 5695
rect 6469 5593 6503 5627
rect 11529 5593 11563 5627
rect 12725 5593 12759 5627
rect 17886 5593 17920 5627
rect 1593 5525 1627 5559
rect 5549 5525 5583 5559
rect 8217 5525 8251 5559
rect 8585 5525 8619 5559
rect 9965 5525 9999 5559
rect 2789 5321 2823 5355
rect 6193 5321 6227 5355
rect 9338 5321 9372 5355
rect 11345 5321 11379 5355
rect 11529 5321 11563 5355
rect 12817 5321 12851 5355
rect 18061 5321 18095 5355
rect 18245 5321 18279 5355
rect 3249 5253 3283 5287
rect 4077 5253 4111 5287
rect 6653 5253 6687 5287
rect 9597 5253 9631 5287
rect 10210 5253 10244 5287
rect 19380 5253 19414 5287
rect 3525 5185 3559 5219
rect 3709 5185 3743 5219
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 8769 5185 8803 5219
rect 8953 5185 8987 5219
rect 9045 5185 9079 5219
rect 9183 5185 9217 5219
rect 9689 5185 9723 5219
rect 11713 5185 11747 5219
rect 11897 5185 11931 5219
rect 20453 5185 20487 5219
rect 4445 5117 4479 5151
rect 4721 5117 4755 5151
rect 6377 5117 6411 5151
rect 9965 5117 9999 5151
rect 12357 5117 12391 5151
rect 12909 5117 12943 5151
rect 13185 5117 13219 5151
rect 14749 5117 14783 5151
rect 15025 5117 15059 5151
rect 19625 5117 19659 5151
rect 2881 5049 2915 5083
rect 4353 5049 4387 5083
rect 8125 5049 8159 5083
rect 12633 5049 12667 5083
rect 14657 5049 14691 5083
rect 3525 4981 3559 5015
rect 16497 4981 16531 5015
rect 20269 4981 20303 5015
rect 6285 4777 6319 4811
rect 9505 4777 9539 4811
rect 13093 4777 13127 4811
rect 13461 4777 13495 4811
rect 14381 4709 14415 4743
rect 5733 4641 5767 4675
rect 4445 4573 4479 4607
rect 4813 4573 4847 4607
rect 6193 4573 6227 4607
rect 8953 4573 8987 4607
rect 9229 4573 9263 4607
rect 9367 4573 9401 4607
rect 12909 4573 12943 4607
rect 13093 4573 13127 4607
rect 13369 4573 13403 4607
rect 4629 4505 4663 4539
rect 4721 4505 4755 4539
rect 5549 4505 5583 4539
rect 9137 4505 9171 4539
rect 14197 4505 14231 4539
rect 4997 4437 5031 4471
rect 7665 4097 7699 4131
rect 7849 4097 7883 4131
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 10057 4097 10091 4131
rect 10154 4097 10188 4131
rect 10701 4097 10735 4131
rect 11713 4097 11747 4131
rect 12541 4097 12575 4131
rect 12725 4097 12759 4131
rect 7941 4029 7975 4063
rect 8217 4029 8251 4063
rect 11989 4029 12023 4063
rect 10333 3961 10367 3995
rect 12357 3961 12391 3995
rect 7665 3893 7699 3927
rect 9689 3893 9723 3927
rect 10609 3893 10643 3927
rect 11621 3893 11655 3927
rect 12449 3893 12483 3927
rect 12541 3893 12575 3927
rect 6009 3689 6043 3723
rect 7192 3689 7226 3723
rect 8677 3689 8711 3723
rect 9965 3689 9999 3723
rect 9505 3621 9539 3655
rect 10149 3553 10183 3587
rect 10425 3553 10459 3587
rect 3985 3485 4019 3519
rect 4077 3485 4111 3519
rect 4261 3485 4295 3519
rect 6929 3485 6963 3519
rect 8953 3485 8987 3519
rect 9367 3485 9401 3519
rect 9781 3485 9815 3519
rect 11989 3485 12023 3519
rect 12245 3485 12279 3519
rect 4537 3417 4571 3451
rect 9137 3417 9171 3451
rect 9229 3417 9263 3451
rect 11897 3349 11931 3383
rect 13369 3349 13403 3383
rect 5273 3145 5307 3179
rect 7849 3145 7883 3179
rect 8953 3145 8987 3179
rect 3801 3077 3835 3111
rect 7757 3009 7791 3043
rect 10701 3009 10735 3043
rect 11800 3009 11834 3043
rect 11897 3009 11931 3043
rect 11989 3009 12023 3043
rect 12173 3009 12207 3043
rect 12357 3009 12391 3043
rect 3525 2941 3559 2975
rect 10425 2941 10459 2975
rect 12633 2941 12667 2975
rect 14197 2941 14231 2975
rect 14473 2941 14507 2975
rect 11621 2873 11655 2907
rect 14105 2873 14139 2907
rect 15945 2805 15979 2839
rect 5457 2601 5491 2635
rect 12633 2601 12667 2635
rect 12909 2601 12943 2635
rect 10701 2465 10735 2499
rect 5273 2397 5307 2431
rect 10425 2397 10459 2431
rect 12449 2397 12483 2431
rect 12817 2397 12851 2431
rect 15761 2397 15795 2431
rect 15577 2329 15611 2363
<< metal1 >>
rect 1104 21786 20792 21808
rect 1104 21734 7214 21786
rect 7266 21734 7278 21786
rect 7330 21734 7342 21786
rect 7394 21734 7406 21786
rect 7458 21734 7470 21786
rect 7522 21734 13214 21786
rect 13266 21734 13278 21786
rect 13330 21734 13342 21786
rect 13394 21734 13406 21786
rect 13458 21734 13470 21786
rect 13522 21734 19214 21786
rect 19266 21734 19278 21786
rect 19330 21734 19342 21786
rect 19394 21734 19406 21786
rect 19458 21734 19470 21786
rect 19522 21734 20792 21786
rect 1104 21712 20792 21734
rect 3326 21496 3332 21548
rect 3384 21496 3390 21548
rect 13814 21496 13820 21548
rect 13872 21536 13878 21548
rect 14093 21539 14151 21545
rect 14093 21536 14105 21539
rect 13872 21508 14105 21536
rect 13872 21496 13878 21508
rect 14093 21505 14105 21508
rect 14139 21505 14151 21539
rect 14093 21499 14151 21505
rect 17770 21496 17776 21548
rect 17828 21496 17834 21548
rect 18049 21539 18107 21545
rect 18049 21505 18061 21539
rect 18095 21536 18107 21539
rect 18138 21536 18144 21548
rect 18095 21508 18144 21536
rect 18095 21505 18107 21508
rect 18049 21499 18107 21505
rect 18138 21496 18144 21508
rect 18196 21496 18202 21548
rect 18690 21496 18696 21548
rect 18748 21536 18754 21548
rect 18969 21539 19027 21545
rect 18969 21536 18981 21539
rect 18748 21508 18981 21536
rect 18748 21496 18754 21508
rect 18969 21505 18981 21508
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 20254 21496 20260 21548
rect 20312 21496 20318 21548
rect 14366 21428 14372 21480
rect 14424 21428 14430 21480
rect 17954 21428 17960 21480
rect 18012 21428 18018 21480
rect 3513 21335 3571 21341
rect 3513 21301 3525 21335
rect 3559 21332 3571 21335
rect 4798 21332 4804 21344
rect 3559 21304 4804 21332
rect 3559 21301 3571 21304
rect 3513 21295 3571 21301
rect 4798 21292 4804 21304
rect 4856 21292 4862 21344
rect 12345 21335 12403 21341
rect 12345 21301 12357 21335
rect 12391 21332 12403 21335
rect 12434 21332 12440 21344
rect 12391 21304 12440 21332
rect 12391 21301 12403 21304
rect 12345 21295 12403 21301
rect 12434 21292 12440 21304
rect 12492 21332 12498 21344
rect 13817 21335 13875 21341
rect 13817 21332 13829 21335
rect 12492 21304 13829 21332
rect 12492 21292 12498 21304
rect 13817 21301 13829 21304
rect 13863 21301 13875 21335
rect 13817 21295 13875 21301
rect 18046 21292 18052 21344
rect 18104 21292 18110 21344
rect 18230 21292 18236 21344
rect 18288 21292 18294 21344
rect 18322 21292 18328 21344
rect 18380 21332 18386 21344
rect 18509 21335 18567 21341
rect 18509 21332 18521 21335
rect 18380 21304 18521 21332
rect 18380 21292 18386 21304
rect 18509 21301 18521 21304
rect 18555 21301 18567 21335
rect 18509 21295 18567 21301
rect 18598 21292 18604 21344
rect 18656 21332 18662 21344
rect 18785 21335 18843 21341
rect 18785 21332 18797 21335
rect 18656 21304 18797 21332
rect 18656 21292 18662 21304
rect 18785 21301 18797 21304
rect 18831 21301 18843 21335
rect 18785 21295 18843 21301
rect 20349 21335 20407 21341
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20438 21332 20444 21344
rect 20395 21304 20444 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 1104 21242 20792 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 10214 21242
rect 10266 21190 10278 21242
rect 10330 21190 10342 21242
rect 10394 21190 10406 21242
rect 10458 21190 10470 21242
rect 10522 21190 16214 21242
rect 16266 21190 16278 21242
rect 16330 21190 16342 21242
rect 16394 21190 16406 21242
rect 16458 21190 16470 21242
rect 16522 21190 20792 21242
rect 1104 21168 20792 21190
rect 12434 21128 12440 21140
rect 12360 21100 12440 21128
rect 5092 20964 8432 20992
rect 5092 20933 5120 20964
rect 8404 20936 8432 20964
rect 5077 20927 5135 20933
rect 5077 20893 5089 20927
rect 5123 20893 5135 20927
rect 5077 20887 5135 20893
rect 6917 20927 6975 20933
rect 6917 20893 6929 20927
rect 6963 20924 6975 20927
rect 7006 20924 7012 20936
rect 6963 20896 7012 20924
rect 6963 20893 6975 20896
rect 6917 20887 6975 20893
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 7098 20884 7104 20936
rect 7156 20884 7162 20936
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 7377 20927 7435 20933
rect 7377 20924 7389 20927
rect 7331 20896 7389 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 7377 20893 7389 20896
rect 7423 20893 7435 20927
rect 7377 20887 7435 20893
rect 8386 20884 8392 20936
rect 8444 20884 8450 20936
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8680 20896 8953 20924
rect 4890 20748 4896 20800
rect 4948 20748 4954 20800
rect 7558 20748 7564 20800
rect 7616 20748 7622 20800
rect 8294 20748 8300 20800
rect 8352 20788 8358 20800
rect 8680 20797 8708 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 12161 20927 12219 20933
rect 12161 20893 12173 20927
rect 12207 20924 12219 20927
rect 12360 20924 12388 21100
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 14366 21088 14372 21140
rect 14424 21088 14430 21140
rect 18046 21088 18052 21140
rect 18104 21128 18110 21140
rect 18693 21131 18751 21137
rect 18693 21128 18705 21131
rect 18104 21100 18705 21128
rect 18104 21088 18110 21100
rect 18693 21097 18705 21100
rect 18739 21128 18751 21131
rect 18782 21128 18788 21140
rect 18739 21100 18788 21128
rect 18739 21097 18751 21100
rect 18693 21091 18751 21097
rect 18782 21088 18788 21100
rect 18840 21088 18846 21140
rect 14384 20992 14412 21088
rect 13832 20964 14412 20992
rect 12618 20924 12624 20936
rect 12207 20896 12624 20924
rect 12207 20893 12219 20896
rect 12161 20887 12219 20893
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 13653 20927 13711 20933
rect 13653 20893 13665 20927
rect 13699 20924 13711 20927
rect 13832 20924 13860 20964
rect 13699 20896 13860 20924
rect 13909 20927 13967 20933
rect 13699 20893 13711 20896
rect 13653 20887 13711 20893
rect 13909 20893 13921 20927
rect 13955 20893 13967 20927
rect 14384 20924 14412 20964
rect 15470 20924 15476 20936
rect 14384 20896 15476 20924
rect 13909 20887 13967 20893
rect 8754 20816 8760 20868
rect 8812 20856 8818 20868
rect 9186 20859 9244 20865
rect 9186 20856 9198 20859
rect 8812 20828 9198 20856
rect 8812 20816 8818 20828
rect 9186 20825 9198 20828
rect 9232 20825 9244 20859
rect 9186 20819 9244 20825
rect 11606 20816 11612 20868
rect 11664 20856 11670 20868
rect 11894 20859 11952 20865
rect 11894 20856 11906 20859
rect 11664 20828 11906 20856
rect 11664 20816 11670 20828
rect 11894 20825 11906 20828
rect 11940 20825 11952 20859
rect 12636 20856 12664 20884
rect 13924 20856 13952 20887
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 15562 20884 15568 20936
rect 15620 20924 15626 20936
rect 17129 20927 17187 20933
rect 17129 20924 17141 20927
rect 15620 20896 17141 20924
rect 15620 20884 15626 20896
rect 17129 20893 17141 20896
rect 17175 20924 17187 20927
rect 17310 20924 17316 20936
rect 17175 20896 17316 20924
rect 17175 20893 17187 20896
rect 17129 20887 17187 20893
rect 17310 20884 17316 20896
rect 17368 20884 17374 20936
rect 12636 20828 13952 20856
rect 11894 20819 11952 20825
rect 15194 20816 15200 20868
rect 15252 20856 15258 20868
rect 15298 20859 15356 20865
rect 15298 20856 15310 20859
rect 15252 20828 15310 20856
rect 15252 20816 15258 20828
rect 15298 20825 15310 20828
rect 15344 20825 15356 20859
rect 15298 20819 15356 20825
rect 17580 20859 17638 20865
rect 17580 20825 17592 20859
rect 17626 20856 17638 20859
rect 17954 20856 17960 20868
rect 17626 20828 17960 20856
rect 17626 20825 17638 20828
rect 17580 20819 17638 20825
rect 17954 20816 17960 20828
rect 18012 20816 18018 20868
rect 8665 20791 8723 20797
rect 8665 20788 8677 20791
rect 8352 20760 8677 20788
rect 8352 20748 8358 20760
rect 8665 20757 8677 20760
rect 8711 20757 8723 20791
rect 8665 20751 8723 20757
rect 10318 20748 10324 20800
rect 10376 20748 10382 20800
rect 10778 20748 10784 20800
rect 10836 20748 10842 20800
rect 12526 20748 12532 20800
rect 12584 20748 12590 20800
rect 14182 20748 14188 20800
rect 14240 20748 14246 20800
rect 1104 20698 20792 20720
rect 1104 20646 7214 20698
rect 7266 20646 7278 20698
rect 7330 20646 7342 20698
rect 7394 20646 7406 20698
rect 7458 20646 7470 20698
rect 7522 20646 13214 20698
rect 13266 20646 13278 20698
rect 13330 20646 13342 20698
rect 13394 20646 13406 20698
rect 13458 20646 13470 20698
rect 13522 20646 19214 20698
rect 19266 20646 19278 20698
rect 19330 20646 19342 20698
rect 19394 20646 19406 20698
rect 19458 20646 19470 20698
rect 19522 20646 20792 20698
rect 1104 20624 20792 20646
rect 8481 20587 8539 20593
rect 8481 20553 8493 20587
rect 8527 20584 8539 20587
rect 8754 20584 8760 20596
rect 8527 20556 8760 20584
rect 8527 20553 8539 20556
rect 8481 20547 8539 20553
rect 8754 20544 8760 20556
rect 8812 20544 8818 20596
rect 11606 20544 11612 20596
rect 11664 20544 11670 20596
rect 6089 20519 6147 20525
rect 6089 20485 6101 20519
rect 6135 20516 6147 20519
rect 6135 20488 7052 20516
rect 6135 20485 6147 20488
rect 6089 20479 6147 20485
rect 7024 20460 7052 20488
rect 7558 20476 7564 20528
rect 7616 20525 7622 20528
rect 7616 20516 7628 20525
rect 7616 20488 7661 20516
rect 7616 20479 7628 20488
rect 7616 20476 7622 20479
rect 10870 20476 10876 20528
rect 10928 20516 10934 20528
rect 11624 20516 11652 20544
rect 12434 20516 12440 20528
rect 10928 20488 12440 20516
rect 10928 20476 10934 20488
rect 12434 20476 12440 20488
rect 12492 20476 12498 20528
rect 12526 20476 12532 20528
rect 12584 20476 12590 20528
rect 12744 20519 12802 20525
rect 12744 20485 12756 20519
rect 12790 20516 12802 20519
rect 14182 20516 14188 20528
rect 12790 20488 14188 20516
rect 12790 20485 12802 20488
rect 12744 20479 12802 20485
rect 14182 20476 14188 20488
rect 14240 20516 14246 20528
rect 16942 20525 16948 20528
rect 14240 20488 14780 20516
rect 14240 20476 14246 20488
rect 4890 20408 4896 20460
rect 4948 20408 4954 20460
rect 5994 20408 6000 20460
rect 6052 20408 6058 20460
rect 6181 20451 6239 20457
rect 6181 20417 6193 20451
rect 6227 20448 6239 20451
rect 6227 20420 6500 20448
rect 6227 20417 6239 20420
rect 6181 20411 6239 20417
rect 4062 20204 4068 20256
rect 4120 20244 4126 20256
rect 4249 20247 4307 20253
rect 4249 20244 4261 20247
rect 4120 20216 4261 20244
rect 4120 20204 4126 20216
rect 4249 20213 4261 20216
rect 4295 20213 4307 20247
rect 4249 20207 4307 20213
rect 5810 20204 5816 20256
rect 5868 20204 5874 20256
rect 6472 20253 6500 20420
rect 7006 20408 7012 20460
rect 7064 20448 7070 20460
rect 8113 20451 8171 20457
rect 7064 20420 8064 20448
rect 7064 20408 7070 20420
rect 8036 20389 8064 20420
rect 8113 20417 8125 20451
rect 8159 20448 8171 20451
rect 8757 20451 8815 20457
rect 8757 20448 8769 20451
rect 8159 20420 8769 20448
rect 8159 20417 8171 20420
rect 8113 20411 8171 20417
rect 8757 20417 8769 20420
rect 8803 20448 8815 20451
rect 10134 20448 10140 20460
rect 8803 20420 10140 20448
rect 8803 20417 8815 20420
rect 8757 20411 8815 20417
rect 10134 20408 10140 20420
rect 10192 20448 10198 20460
rect 10318 20448 10324 20460
rect 10192 20420 10324 20448
rect 10192 20408 10198 20420
rect 10318 20408 10324 20420
rect 10376 20448 10382 20460
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10376 20420 10517 20448
rect 10376 20408 10382 20420
rect 10505 20417 10517 20420
rect 10551 20448 10563 20451
rect 11241 20451 11299 20457
rect 11241 20448 11253 20451
rect 10551 20420 11253 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 11241 20417 11253 20420
rect 11287 20448 11299 20451
rect 12544 20448 12572 20476
rect 13337 20451 13395 20457
rect 13337 20448 13349 20451
rect 11287 20420 12020 20448
rect 12544 20420 13349 20448
rect 11287 20417 11299 20420
rect 11241 20411 11299 20417
rect 7837 20383 7895 20389
rect 7837 20349 7849 20383
rect 7883 20349 7895 20383
rect 7837 20343 7895 20349
rect 8021 20383 8079 20389
rect 8021 20349 8033 20383
rect 8067 20349 8079 20383
rect 8021 20343 8079 20349
rect 7852 20312 7880 20343
rect 8294 20340 8300 20392
rect 8352 20340 8358 20392
rect 8312 20312 8340 20340
rect 7852 20284 8340 20312
rect 6457 20247 6515 20253
rect 6457 20213 6469 20247
rect 6503 20244 6515 20247
rect 6546 20244 6552 20256
rect 6503 20216 6552 20244
rect 6503 20213 6515 20216
rect 6457 20207 6515 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 11992 20244 12020 20420
rect 13337 20417 13349 20420
rect 13383 20448 13395 20451
rect 13722 20448 13728 20460
rect 13383 20420 13728 20448
rect 13383 20417 13395 20420
rect 13337 20411 13395 20417
rect 13722 20408 13728 20420
rect 13780 20448 13786 20460
rect 14752 20457 14780 20488
rect 16936 20479 16948 20525
rect 17000 20516 17006 20528
rect 17770 20516 17776 20528
rect 17000 20488 17776 20516
rect 16942 20476 16948 20479
rect 17000 20476 17006 20488
rect 17770 20476 17776 20488
rect 17828 20476 17834 20528
rect 18138 20476 18144 20528
rect 18196 20516 18202 20528
rect 18478 20519 18536 20525
rect 18478 20516 18490 20519
rect 18196 20488 18490 20516
rect 18196 20476 18202 20488
rect 18478 20485 18490 20488
rect 18524 20485 18536 20519
rect 18478 20479 18536 20485
rect 14645 20451 14703 20457
rect 14645 20448 14657 20451
rect 13780 20420 14657 20448
rect 13780 20408 13786 20420
rect 14645 20417 14657 20420
rect 14691 20417 14703 20451
rect 14645 20411 14703 20417
rect 14737 20451 14795 20457
rect 14737 20417 14749 20451
rect 14783 20417 14795 20451
rect 14737 20411 14795 20417
rect 17310 20408 17316 20460
rect 17368 20448 17374 20460
rect 18233 20451 18291 20457
rect 18233 20448 18245 20451
rect 17368 20420 18245 20448
rect 17368 20408 17374 20420
rect 18233 20417 18245 20420
rect 18279 20448 18291 20451
rect 18322 20448 18328 20460
rect 18279 20420 18328 20448
rect 18279 20417 18291 20420
rect 18233 20411 18291 20417
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 13035 20352 13093 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 16669 20383 16727 20389
rect 16669 20380 16681 20383
rect 13081 20343 13139 20349
rect 16408 20352 16681 20380
rect 12618 20244 12624 20256
rect 11992 20216 12624 20244
rect 12618 20204 12624 20216
rect 12676 20244 12682 20256
rect 13004 20244 13032 20343
rect 14461 20315 14519 20321
rect 14461 20281 14473 20315
rect 14507 20312 14519 20315
rect 14507 20284 15240 20312
rect 14507 20281 14519 20284
rect 14461 20275 14519 20281
rect 14844 20253 14872 20284
rect 15212 20256 15240 20284
rect 12676 20216 13032 20244
rect 14829 20247 14887 20253
rect 12676 20204 12682 20216
rect 14829 20213 14841 20247
rect 14875 20213 14887 20247
rect 14829 20207 14887 20213
rect 15010 20204 15016 20256
rect 15068 20204 15074 20256
rect 15194 20204 15200 20256
rect 15252 20204 15258 20256
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 16408 20253 16436 20352
rect 16669 20349 16681 20352
rect 16715 20349 16727 20383
rect 16669 20343 16727 20349
rect 16393 20247 16451 20253
rect 16393 20244 16405 20247
rect 15620 20216 16405 20244
rect 15620 20204 15626 20216
rect 16393 20213 16405 20216
rect 16439 20213 16451 20247
rect 16393 20207 16451 20213
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 18049 20247 18107 20253
rect 18049 20244 18061 20247
rect 18012 20216 18061 20244
rect 18012 20204 18018 20216
rect 18049 20213 18061 20216
rect 18095 20213 18107 20247
rect 18049 20207 18107 20213
rect 19610 20204 19616 20256
rect 19668 20204 19674 20256
rect 1104 20154 20792 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 10214 20154
rect 10266 20102 10278 20154
rect 10330 20102 10342 20154
rect 10394 20102 10406 20154
rect 10458 20102 10470 20154
rect 10522 20102 16214 20154
rect 16266 20102 16278 20154
rect 16330 20102 16342 20154
rect 16394 20102 16406 20154
rect 16458 20102 16470 20154
rect 16522 20102 20792 20154
rect 1104 20080 20792 20102
rect 7098 20000 7104 20052
rect 7156 20040 7162 20052
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 7156 20012 7297 20040
rect 7156 20000 7162 20012
rect 7285 20009 7297 20012
rect 7331 20009 7343 20043
rect 7285 20003 7343 20009
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 10192 20012 10333 20040
rect 10192 20000 10198 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 10321 20003 10379 20009
rect 10336 19904 10364 20003
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 12894 20040 12900 20052
rect 12676 20012 12900 20040
rect 12676 20000 12682 20012
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 14277 20043 14335 20049
rect 14277 20009 14289 20043
rect 14323 20040 14335 20043
rect 15194 20040 15200 20052
rect 14323 20012 15200 20040
rect 14323 20009 14335 20012
rect 14277 20003 14335 20009
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 16942 20000 16948 20052
rect 17000 20000 17006 20052
rect 17310 20000 17316 20052
rect 17368 20040 17374 20052
rect 17405 20043 17463 20049
rect 17405 20040 17417 20043
rect 17368 20012 17417 20040
rect 17368 20000 17374 20012
rect 17405 20009 17417 20012
rect 17451 20009 17463 20043
rect 17405 20003 17463 20009
rect 17681 20043 17739 20049
rect 17681 20009 17693 20043
rect 17727 20040 17739 20043
rect 18138 20040 18144 20052
rect 17727 20012 18144 20040
rect 17727 20009 17739 20012
rect 17681 20003 17739 20009
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 18322 20000 18328 20052
rect 18380 20040 18386 20052
rect 18380 20012 19104 20040
rect 18380 20000 18386 20012
rect 19076 19913 19104 20012
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 10336 19876 10517 19904
rect 10505 19873 10517 19876
rect 10551 19873 10563 19907
rect 10505 19867 10563 19873
rect 19061 19907 19119 19913
rect 19061 19873 19073 19907
rect 19107 19873 19119 19907
rect 19061 19867 19119 19873
rect 4062 19796 4068 19848
rect 4120 19796 4126 19848
rect 5994 19796 6000 19848
rect 6052 19796 6058 19848
rect 6270 19796 6276 19848
rect 6328 19796 6334 19848
rect 6454 19836 6460 19848
rect 6380 19808 6460 19836
rect 6012 19768 6040 19796
rect 6380 19768 6408 19808
rect 6454 19796 6460 19808
rect 6512 19796 6518 19848
rect 6546 19796 6552 19848
rect 6604 19836 6610 19848
rect 10778 19845 10784 19848
rect 7101 19839 7159 19845
rect 7101 19836 7113 19839
rect 6604 19808 7113 19836
rect 6604 19796 6610 19808
rect 7101 19805 7113 19808
rect 7147 19805 7159 19839
rect 10772 19836 10784 19845
rect 10739 19808 10784 19836
rect 7101 19799 7159 19805
rect 10772 19799 10784 19808
rect 10836 19836 10842 19848
rect 10836 19808 12204 19836
rect 10778 19796 10784 19799
rect 10836 19796 10842 19808
rect 6917 19771 6975 19777
rect 6917 19768 6929 19771
rect 6012 19740 6929 19768
rect 6917 19737 6929 19740
rect 6963 19737 6975 19771
rect 6917 19731 6975 19737
rect 11790 19728 11796 19780
rect 11848 19768 11854 19780
rect 12069 19771 12127 19777
rect 12069 19768 12081 19771
rect 11848 19740 12081 19768
rect 11848 19728 11854 19740
rect 12069 19737 12081 19740
rect 12115 19737 12127 19771
rect 12176 19768 12204 19808
rect 12434 19796 12440 19848
rect 12492 19796 12498 19848
rect 13722 19796 13728 19848
rect 13780 19836 13786 19848
rect 13780 19808 13952 19836
rect 13780 19796 13786 19808
rect 12345 19771 12403 19777
rect 12345 19768 12357 19771
rect 12176 19740 12357 19768
rect 12069 19731 12127 19737
rect 12345 19737 12357 19740
rect 12391 19737 12403 19771
rect 12345 19731 12403 19737
rect 4062 19660 4068 19712
rect 4120 19660 4126 19712
rect 6362 19660 6368 19712
rect 6420 19660 6426 19712
rect 11146 19660 11152 19712
rect 11204 19700 11210 19712
rect 11885 19703 11943 19709
rect 11885 19700 11897 19703
rect 11204 19672 11897 19700
rect 11204 19660 11210 19672
rect 11885 19669 11897 19672
rect 11931 19700 11943 19703
rect 12250 19700 12256 19712
rect 11931 19672 12256 19700
rect 11931 19669 11943 19672
rect 11885 19663 11943 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12452 19709 12480 19796
rect 12621 19771 12679 19777
rect 12621 19737 12633 19771
rect 12667 19768 12679 19771
rect 13814 19768 13820 19780
rect 12667 19740 13820 19768
rect 12667 19737 12679 19740
rect 12621 19731 12679 19737
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 13924 19768 13952 19808
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 15562 19836 15568 19848
rect 14240 19808 14504 19836
rect 14240 19796 14246 19808
rect 14476 19777 14504 19808
rect 15396 19808 15568 19836
rect 14461 19771 14519 19777
rect 13924 19740 14228 19768
rect 12437 19703 12495 19709
rect 12437 19669 12449 19703
rect 12483 19669 12495 19703
rect 12437 19663 12495 19669
rect 14090 19660 14096 19712
rect 14148 19660 14154 19712
rect 14200 19700 14228 19740
rect 14461 19737 14473 19771
rect 14507 19737 14519 19771
rect 14461 19731 14519 19737
rect 15396 19712 15424 19808
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 18782 19796 18788 19848
rect 18840 19845 18846 19848
rect 18840 19836 18852 19845
rect 18840 19808 18885 19836
rect 18840 19799 18852 19808
rect 18840 19796 18846 19799
rect 15832 19771 15890 19777
rect 15832 19737 15844 19771
rect 15878 19768 15890 19771
rect 16114 19768 16120 19780
rect 15878 19740 16120 19768
rect 15878 19737 15890 19740
rect 15832 19731 15890 19737
rect 16114 19728 16120 19740
rect 16172 19728 16178 19780
rect 14256 19703 14314 19709
rect 14256 19700 14268 19703
rect 14200 19672 14268 19700
rect 14256 19669 14268 19672
rect 14302 19669 14314 19703
rect 14256 19663 14314 19669
rect 15378 19660 15384 19712
rect 15436 19660 15442 19712
rect 1104 19610 20792 19632
rect 1104 19558 7214 19610
rect 7266 19558 7278 19610
rect 7330 19558 7342 19610
rect 7394 19558 7406 19610
rect 7458 19558 7470 19610
rect 7522 19558 13214 19610
rect 13266 19558 13278 19610
rect 13330 19558 13342 19610
rect 13394 19558 13406 19610
rect 13458 19558 13470 19610
rect 13522 19558 19214 19610
rect 19266 19558 19278 19610
rect 19330 19558 19342 19610
rect 19394 19558 19406 19610
rect 19458 19558 19470 19610
rect 19522 19558 20792 19610
rect 1104 19536 20792 19558
rect 4062 19496 4068 19508
rect 2746 19468 4068 19496
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 2746 19360 2774 19468
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 6082 19499 6140 19505
rect 6082 19465 6094 19499
rect 6128 19496 6140 19499
rect 6270 19496 6276 19508
rect 6128 19468 6276 19496
rect 6128 19465 6140 19468
rect 6082 19459 6140 19465
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 6362 19456 6368 19508
rect 6420 19456 6426 19508
rect 9306 19456 9312 19508
rect 9364 19496 9370 19508
rect 10045 19499 10103 19505
rect 10045 19496 10057 19499
rect 9364 19468 10057 19496
rect 9364 19456 9370 19468
rect 10045 19465 10057 19468
rect 10091 19465 10103 19499
rect 10045 19459 10103 19465
rect 11333 19499 11391 19505
rect 11333 19465 11345 19499
rect 11379 19496 11391 19499
rect 11379 19468 13584 19496
rect 11379 19465 11391 19468
rect 11333 19459 11391 19465
rect 6380 19428 6408 19456
rect 7570 19431 7628 19437
rect 7570 19428 7582 19431
rect 6380 19400 7582 19428
rect 7570 19397 7582 19400
rect 7616 19397 7628 19431
rect 7570 19391 7628 19397
rect 10796 19400 11100 19428
rect 10796 19372 10824 19400
rect 4614 19369 4620 19372
rect 2547 19332 2774 19360
rect 3145 19363 3203 19369
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 3145 19329 3157 19363
rect 3191 19360 3203 19363
rect 3237 19363 3295 19369
rect 3237 19360 3249 19363
rect 3191 19332 3249 19360
rect 3191 19329 3203 19332
rect 3145 19323 3203 19329
rect 3237 19329 3249 19332
rect 3283 19329 3295 19363
rect 3237 19323 3295 19329
rect 4608 19323 4620 19369
rect 4614 19320 4620 19323
rect 4672 19320 4678 19372
rect 5902 19320 5908 19372
rect 5960 19320 5966 19372
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19329 6055 19363
rect 5997 19323 6055 19329
rect 6181 19363 6239 19369
rect 6181 19329 6193 19363
rect 6227 19360 6239 19363
rect 6270 19360 6276 19372
rect 6227 19332 6276 19360
rect 6227 19329 6239 19332
rect 6181 19323 6239 19329
rect 4341 19295 4399 19301
rect 4341 19292 4353 19295
rect 4172 19264 4353 19292
rect 3234 19116 3240 19168
rect 3292 19116 3298 19168
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4172 19165 4200 19264
rect 4341 19261 4353 19264
rect 4387 19261 4399 19295
rect 6012 19292 6040 19323
rect 6270 19320 6276 19332
rect 6328 19360 6334 19372
rect 8294 19360 8300 19372
rect 6328 19332 6500 19360
rect 6328 19320 6334 19332
rect 4341 19255 4399 19261
rect 5736 19264 6040 19292
rect 5736 19168 5764 19264
rect 6472 19233 6500 19332
rect 8220 19332 8300 19360
rect 7837 19295 7895 19301
rect 7837 19261 7849 19295
rect 7883 19292 7895 19295
rect 8113 19295 8171 19301
rect 8113 19292 8125 19295
rect 7883 19264 8125 19292
rect 7883 19261 7895 19264
rect 7837 19255 7895 19261
rect 8113 19261 8125 19264
rect 8159 19292 8171 19295
rect 8220 19292 8248 19332
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 10042 19360 10048 19372
rect 9706 19332 10048 19360
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 10778 19320 10784 19372
rect 10836 19320 10842 19372
rect 10870 19320 10876 19372
rect 10928 19320 10934 19372
rect 11072 19369 11100 19400
rect 12250 19388 12256 19440
rect 12308 19428 12314 19440
rect 12722 19431 12780 19437
rect 12722 19428 12734 19431
rect 12308 19400 12734 19428
rect 12308 19388 12314 19400
rect 12722 19397 12734 19400
rect 12768 19397 12780 19431
rect 12722 19391 12780 19397
rect 12894 19388 12900 19440
rect 12952 19388 12958 19440
rect 11057 19363 11115 19369
rect 11057 19329 11069 19363
rect 11103 19329 11115 19363
rect 11057 19323 11115 19329
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 12912 19360 12940 19388
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 11195 19332 11836 19360
rect 12912 19332 13001 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 8159 19264 8248 19292
rect 8159 19261 8171 19264
rect 8113 19255 8171 19261
rect 6457 19227 6515 19233
rect 6457 19193 6469 19227
rect 6503 19193 6515 19227
rect 6457 19187 6515 19193
rect 7852 19168 7880 19255
rect 8570 19252 8576 19304
rect 8628 19252 8634 19304
rect 11808 19236 11836 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 13556 19360 13584 19468
rect 14090 19456 14096 19508
rect 14148 19456 14154 19508
rect 15013 19499 15071 19505
rect 15013 19465 15025 19499
rect 15059 19496 15071 19499
rect 15562 19496 15568 19508
rect 15059 19468 15568 19496
rect 15059 19465 15071 19468
rect 15013 19459 15071 19465
rect 15562 19456 15568 19468
rect 15620 19456 15626 19508
rect 17770 19456 17776 19508
rect 17828 19496 17834 19508
rect 17865 19499 17923 19505
rect 17865 19496 17877 19499
rect 17828 19468 17877 19496
rect 17828 19456 17834 19468
rect 17865 19465 17877 19468
rect 17911 19465 17923 19499
rect 17865 19459 17923 19465
rect 17954 19456 17960 19508
rect 18012 19456 18018 19508
rect 18049 19499 18107 19505
rect 18049 19465 18061 19499
rect 18095 19496 18107 19499
rect 18782 19496 18788 19508
rect 18095 19468 18788 19496
rect 18095 19465 18107 19468
rect 18049 19459 18107 19465
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 14108 19428 14136 19456
rect 14185 19431 14243 19437
rect 14185 19428 14197 19431
rect 14108 19400 14197 19428
rect 14185 19397 14197 19400
rect 14231 19397 14243 19431
rect 14185 19391 14243 19397
rect 14401 19431 14459 19437
rect 14401 19397 14413 19431
rect 14447 19428 14459 19431
rect 14550 19428 14556 19440
rect 14447 19400 14556 19428
rect 14447 19397 14459 19400
rect 14401 19391 14459 19397
rect 14550 19388 14556 19400
rect 14608 19388 14614 19440
rect 15930 19428 15936 19440
rect 14660 19400 15936 19428
rect 14660 19369 14688 19400
rect 15930 19388 15936 19400
rect 15988 19388 15994 19440
rect 18138 19388 18144 19440
rect 18196 19428 18202 19440
rect 18233 19431 18291 19437
rect 18233 19428 18245 19431
rect 18196 19400 18245 19428
rect 18196 19388 18202 19400
rect 18233 19397 18245 19400
rect 18279 19397 18291 19431
rect 18233 19391 18291 19397
rect 18322 19388 18328 19440
rect 18380 19428 18386 19440
rect 18877 19431 18935 19437
rect 18877 19428 18889 19431
rect 18380 19400 18889 19428
rect 18380 19388 18386 19400
rect 18877 19397 18889 19400
rect 18923 19397 18935 19431
rect 18877 19391 18935 19397
rect 14645 19363 14703 19369
rect 13556 19332 14504 19360
rect 12989 19323 13047 19329
rect 11790 19184 11796 19236
rect 11848 19184 11854 19236
rect 4157 19159 4215 19165
rect 4157 19156 4169 19159
rect 4120 19128 4169 19156
rect 4120 19116 4126 19128
rect 4157 19125 4169 19128
rect 4203 19125 4215 19159
rect 4157 19119 4215 19125
rect 5718 19116 5724 19168
rect 5776 19116 5782 19168
rect 7834 19116 7840 19168
rect 7892 19116 7898 19168
rect 10778 19116 10784 19168
rect 10836 19116 10842 19168
rect 11146 19116 11152 19168
rect 11204 19116 11210 19168
rect 11609 19159 11667 19165
rect 11609 19125 11621 19159
rect 11655 19156 11667 19159
rect 11808 19156 11836 19184
rect 11655 19128 11836 19156
rect 11655 19125 11667 19128
rect 11609 19119 11667 19125
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14369 19159 14427 19165
rect 14369 19156 14381 19159
rect 13872 19128 14381 19156
rect 13872 19116 13878 19128
rect 14369 19125 14381 19128
rect 14415 19125 14427 19159
rect 14476 19156 14504 19332
rect 14645 19329 14657 19363
rect 14691 19329 14703 19363
rect 14645 19323 14703 19329
rect 14829 19363 14887 19369
rect 14829 19329 14841 19363
rect 14875 19360 14887 19363
rect 15010 19360 15016 19372
rect 14875 19332 15016 19360
rect 14875 19329 14887 19332
rect 14829 19323 14887 19329
rect 15010 19320 15016 19332
rect 15068 19320 15074 19372
rect 18892 19360 18920 19391
rect 19610 19388 19616 19440
rect 19668 19428 19674 19440
rect 20174 19431 20232 19437
rect 20174 19428 20186 19431
rect 19668 19400 20186 19428
rect 19668 19388 19674 19400
rect 20174 19397 20186 19400
rect 20220 19397 20232 19431
rect 20174 19391 20232 19397
rect 20441 19363 20499 19369
rect 20441 19360 20453 19363
rect 18892 19332 20453 19360
rect 20441 19329 20453 19332
rect 20487 19329 20499 19363
rect 20441 19323 20499 19329
rect 14553 19227 14611 19233
rect 14553 19193 14565 19227
rect 14599 19224 14611 19227
rect 15194 19224 15200 19236
rect 14599 19196 15200 19224
rect 14599 19193 14611 19196
rect 14553 19187 14611 19193
rect 15194 19184 15200 19196
rect 15252 19184 15258 19236
rect 14645 19159 14703 19165
rect 14645 19156 14657 19159
rect 14476 19128 14657 19156
rect 14369 19119 14427 19125
rect 14645 19125 14657 19128
rect 14691 19125 14703 19159
rect 14645 19119 14703 19125
rect 17681 19159 17739 19165
rect 17681 19125 17693 19159
rect 17727 19156 17739 19159
rect 17954 19156 17960 19168
rect 17727 19128 17960 19156
rect 17727 19125 17739 19128
rect 17681 19119 17739 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 19061 19159 19119 19165
rect 19061 19125 19073 19159
rect 19107 19156 19119 19159
rect 19794 19156 19800 19168
rect 19107 19128 19800 19156
rect 19107 19125 19119 19128
rect 19061 19119 19119 19125
rect 19794 19116 19800 19128
rect 19852 19116 19858 19168
rect 1104 19066 20792 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 10214 19066
rect 10266 19014 10278 19066
rect 10330 19014 10342 19066
rect 10394 19014 10406 19066
rect 10458 19014 10470 19066
rect 10522 19014 16214 19066
rect 16266 19014 16278 19066
rect 16330 19014 16342 19066
rect 16394 19014 16406 19066
rect 16458 19014 16470 19066
rect 16522 19014 20792 19066
rect 1104 18992 20792 19014
rect 3234 18952 3240 18964
rect 2746 18924 3240 18952
rect 2746 18816 2774 18924
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 4154 18912 4160 18964
rect 4212 18912 4218 18964
rect 4525 18955 4583 18961
rect 4525 18921 4537 18955
rect 4571 18952 4583 18955
rect 4614 18952 4620 18964
rect 4571 18924 4620 18952
rect 4571 18921 4583 18924
rect 4525 18915 4583 18921
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 6270 18912 6276 18964
rect 6328 18912 6334 18964
rect 6454 18912 6460 18964
rect 6512 18912 6518 18964
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 9033 18955 9091 18961
rect 9033 18952 9045 18955
rect 8628 18924 9045 18952
rect 8628 18912 8634 18924
rect 9033 18921 9045 18924
rect 9079 18921 9091 18955
rect 9033 18915 9091 18921
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 11241 18955 11299 18961
rect 11241 18952 11253 18955
rect 10836 18924 11253 18952
rect 10836 18912 10842 18924
rect 11241 18921 11253 18924
rect 11287 18952 11299 18955
rect 12434 18952 12440 18964
rect 11287 18924 12440 18952
rect 11287 18921 11299 18924
rect 11241 18915 11299 18921
rect 4172 18884 4200 18912
rect 5810 18884 5816 18896
rect 4172 18856 5816 18884
rect 5810 18844 5816 18856
rect 5868 18884 5874 18896
rect 6733 18887 6791 18893
rect 6733 18884 6745 18887
rect 5868 18856 6745 18884
rect 5868 18844 5874 18856
rect 6733 18853 6745 18856
rect 6779 18884 6791 18887
rect 7834 18884 7840 18896
rect 6779 18856 7840 18884
rect 6779 18853 6791 18856
rect 6733 18847 6791 18853
rect 7834 18844 7840 18856
rect 7892 18844 7898 18896
rect 1964 18788 2774 18816
rect 4985 18819 5043 18825
rect 1964 18757 1992 18788
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 5166 18816 5172 18828
rect 5031 18788 5172 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 5166 18776 5172 18788
rect 5224 18816 5230 18828
rect 5902 18816 5908 18828
rect 5224 18788 5908 18816
rect 5224 18776 5230 18788
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 9306 18776 9312 18828
rect 9364 18776 9370 18828
rect 11256 18816 11284 18915
rect 12434 18912 12440 18924
rect 12492 18952 12498 18964
rect 12894 18952 12900 18964
rect 12492 18924 12900 18952
rect 12492 18912 12498 18924
rect 12894 18912 12900 18924
rect 12952 18952 12958 18964
rect 13722 18952 13728 18964
rect 12952 18924 13728 18952
rect 12952 18912 12958 18924
rect 13722 18912 13728 18924
rect 13780 18952 13786 18964
rect 13817 18955 13875 18961
rect 13817 18952 13829 18955
rect 13780 18924 13829 18952
rect 13780 18912 13786 18924
rect 13817 18921 13829 18924
rect 13863 18952 13875 18955
rect 15289 18955 15347 18961
rect 15289 18952 15301 18955
rect 13863 18924 15301 18952
rect 13863 18921 13875 18924
rect 13817 18915 13875 18921
rect 15289 18921 15301 18924
rect 15335 18921 15347 18955
rect 15289 18915 15347 18921
rect 12805 18887 12863 18893
rect 12805 18853 12817 18887
rect 12851 18884 12863 18887
rect 12851 18856 14228 18884
rect 12851 18853 12863 18856
rect 12805 18847 12863 18853
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11256 18788 11437 18816
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 1949 18751 2007 18757
rect 1949 18717 1961 18751
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18748 2651 18751
rect 2685 18751 2743 18757
rect 2685 18748 2697 18751
rect 2639 18720 2697 18748
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 2685 18717 2697 18720
rect 2731 18717 2743 18751
rect 2685 18711 2743 18717
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18748 4951 18751
rect 5718 18748 5724 18760
rect 4939 18720 5724 18748
rect 4939 18717 4951 18720
rect 4893 18711 4951 18717
rect 5718 18708 5724 18720
rect 5776 18748 5782 18760
rect 9125 18751 9183 18757
rect 5776 18720 6132 18748
rect 5776 18708 5782 18720
rect 5902 18640 5908 18692
rect 5960 18640 5966 18692
rect 6104 18689 6132 18720
rect 9125 18717 9137 18751
rect 9171 18748 9183 18751
rect 9324 18748 9352 18776
rect 9171 18720 9352 18748
rect 9171 18717 9183 18720
rect 9125 18711 9183 18717
rect 6089 18683 6147 18689
rect 6089 18649 6101 18683
rect 6135 18649 6147 18683
rect 6089 18643 6147 18649
rect 11692 18683 11750 18689
rect 11692 18649 11704 18683
rect 11738 18680 11750 18683
rect 11790 18680 11796 18692
rect 11738 18652 11796 18680
rect 11738 18649 11750 18652
rect 11692 18643 11750 18649
rect 11790 18640 11796 18652
rect 11848 18640 11854 18692
rect 14090 18640 14096 18692
rect 14148 18640 14154 18692
rect 14200 18680 14228 18856
rect 14550 18844 14556 18896
rect 14608 18884 14614 18896
rect 14608 18856 14688 18884
rect 14608 18844 14614 18856
rect 14660 18825 14688 18856
rect 14645 18819 14703 18825
rect 14645 18785 14657 18819
rect 14691 18785 14703 18819
rect 15304 18816 15332 18915
rect 16942 18912 16948 18964
rect 17000 18912 17006 18964
rect 18230 18912 18236 18964
rect 18288 18952 18294 18964
rect 18325 18955 18383 18961
rect 18325 18952 18337 18955
rect 18288 18924 18337 18952
rect 18288 18912 18294 18924
rect 18325 18921 18337 18924
rect 18371 18921 18383 18955
rect 18325 18915 18383 18921
rect 19610 18912 19616 18964
rect 19668 18912 19674 18964
rect 17313 18887 17371 18893
rect 17313 18853 17325 18887
rect 17359 18853 17371 18887
rect 17313 18847 17371 18853
rect 15378 18816 15384 18828
rect 15304 18788 15384 18816
rect 14645 18779 14703 18785
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 17037 18819 17095 18825
rect 17037 18816 17049 18819
rect 16408 18788 17049 18816
rect 15470 18708 15476 18760
rect 15528 18748 15534 18760
rect 15637 18751 15695 18757
rect 15637 18748 15649 18751
rect 15528 18720 15649 18748
rect 15528 18708 15534 18720
rect 15637 18717 15649 18720
rect 15683 18717 15695 18751
rect 15637 18711 15695 18717
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 16408 18748 16436 18788
rect 17037 18785 17049 18788
rect 17083 18785 17095 18819
rect 17328 18816 17356 18847
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 17328 18788 18429 18816
rect 17037 18779 17095 18785
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 19613 18819 19671 18825
rect 19613 18785 19625 18819
rect 19659 18816 19671 18819
rect 19659 18788 19840 18816
rect 19659 18785 19671 18788
rect 19613 18779 19671 18785
rect 19812 18760 19840 18788
rect 16172 18720 16436 18748
rect 16945 18751 17003 18757
rect 16172 18708 16178 18720
rect 16945 18717 16957 18751
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 19429 18751 19487 18757
rect 18555 18720 19288 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 16960 18680 16988 18711
rect 14200 18652 14504 18680
rect 16960 18652 17080 18680
rect 2866 18572 2872 18624
rect 2924 18572 2930 18624
rect 5920 18612 5948 18640
rect 14476 18624 14504 18652
rect 17052 18624 17080 18652
rect 6289 18615 6347 18621
rect 6289 18612 6301 18615
rect 5920 18584 6301 18612
rect 6289 18581 6301 18584
rect 6335 18581 6347 18615
rect 6289 18575 6347 18581
rect 14182 18572 14188 18624
rect 14240 18612 14246 18624
rect 14277 18615 14335 18621
rect 14277 18612 14289 18615
rect 14240 18584 14289 18612
rect 14240 18572 14246 18584
rect 14277 18581 14289 18584
rect 14323 18581 14335 18615
rect 14277 18575 14335 18581
rect 14366 18572 14372 18624
rect 14424 18572 14430 18624
rect 14458 18572 14464 18624
rect 14516 18572 14522 18624
rect 16761 18615 16819 18621
rect 16761 18581 16773 18615
rect 16807 18612 16819 18615
rect 17034 18612 17040 18624
rect 16807 18584 17040 18612
rect 16807 18581 16819 18584
rect 16761 18575 16819 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 18138 18572 18144 18624
rect 18196 18572 18202 18624
rect 19260 18621 19288 18720
rect 19429 18717 19441 18751
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 19444 18680 19472 18711
rect 19702 18708 19708 18760
rect 19760 18708 19766 18760
rect 19794 18708 19800 18760
rect 19852 18708 19858 18760
rect 19886 18708 19892 18760
rect 19944 18708 19950 18760
rect 19904 18680 19932 18708
rect 19444 18652 19932 18680
rect 19245 18615 19303 18621
rect 19245 18581 19257 18615
rect 19291 18581 19303 18615
rect 19245 18575 19303 18581
rect 1104 18522 20792 18544
rect 1104 18470 7214 18522
rect 7266 18470 7278 18522
rect 7330 18470 7342 18522
rect 7394 18470 7406 18522
rect 7458 18470 7470 18522
rect 7522 18470 13214 18522
rect 13266 18470 13278 18522
rect 13330 18470 13342 18522
rect 13394 18470 13406 18522
rect 13458 18470 13470 18522
rect 13522 18470 19214 18522
rect 19266 18470 19278 18522
rect 19330 18470 19342 18522
rect 19394 18470 19406 18522
rect 19458 18470 19470 18522
rect 19522 18470 20792 18522
rect 1104 18448 20792 18470
rect 9306 18408 9312 18420
rect 7668 18380 9312 18408
rect 7561 18275 7619 18281
rect 7561 18241 7573 18275
rect 7607 18241 7619 18275
rect 7561 18235 7619 18241
rect 4706 18164 4712 18216
rect 4764 18164 4770 18216
rect 7576 18068 7604 18235
rect 7668 18213 7696 18380
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 12253 18411 12311 18417
rect 12253 18377 12265 18411
rect 12299 18408 12311 18411
rect 12434 18408 12440 18420
rect 12299 18380 12440 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 8018 18232 8024 18284
rect 8076 18232 8082 18284
rect 10042 18272 10048 18284
rect 9430 18244 10048 18272
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 12360 18281 12388 18380
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 14366 18408 14372 18420
rect 13771 18380 14372 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 14700 18380 15792 18408
rect 14700 18368 14706 18380
rect 12612 18343 12670 18349
rect 12612 18309 12624 18343
rect 12658 18340 12670 18343
rect 14458 18340 14464 18352
rect 12658 18312 14464 18340
rect 12658 18309 12670 18312
rect 12612 18303 12670 18309
rect 14458 18300 14464 18312
rect 14516 18340 14522 18352
rect 15473 18343 15531 18349
rect 15473 18340 15485 18343
rect 14516 18312 15485 18340
rect 14516 18300 14522 18312
rect 15473 18309 15485 18312
rect 15519 18309 15531 18343
rect 15473 18303 15531 18309
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 15764 18281 15792 18380
rect 15930 18368 15936 18420
rect 15988 18368 15994 18420
rect 16761 18411 16819 18417
rect 16761 18377 16773 18411
rect 16807 18408 16819 18411
rect 16942 18408 16948 18420
rect 16807 18380 16948 18408
rect 16807 18377 16819 18380
rect 16761 18371 16819 18377
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 19610 18368 19616 18420
rect 19668 18368 19674 18420
rect 16114 18300 16120 18352
rect 16172 18300 16178 18352
rect 16333 18343 16391 18349
rect 16333 18309 16345 18343
rect 16379 18340 16391 18343
rect 17034 18340 17040 18352
rect 16379 18312 17040 18340
rect 16379 18309 16391 18312
rect 16333 18303 16391 18309
rect 17034 18300 17040 18312
rect 17092 18340 17098 18352
rect 17874 18343 17932 18349
rect 17874 18340 17886 18343
rect 17092 18312 17886 18340
rect 17092 18300 17098 18312
rect 17874 18309 17886 18312
rect 17920 18309 17932 18343
rect 17874 18303 17932 18309
rect 18500 18343 18558 18349
rect 18500 18309 18512 18343
rect 18546 18340 18558 18343
rect 19794 18340 19800 18352
rect 18546 18312 19800 18340
rect 18546 18309 18558 18312
rect 18500 18303 18558 18309
rect 19794 18300 19800 18312
rect 19852 18300 19858 18352
rect 15114 18275 15172 18281
rect 15114 18272 15126 18275
rect 14240 18244 15126 18272
rect 14240 18232 14246 18244
rect 15114 18241 15126 18244
rect 15160 18272 15172 18275
rect 15749 18275 15807 18281
rect 15160 18244 15516 18272
rect 15160 18241 15172 18244
rect 15114 18235 15172 18241
rect 7653 18207 7711 18213
rect 7653 18173 7665 18207
rect 7699 18173 7711 18207
rect 8297 18207 8355 18213
rect 8297 18204 8309 18207
rect 7653 18167 7711 18173
rect 8128 18176 8309 18204
rect 7929 18139 7987 18145
rect 7929 18105 7941 18139
rect 7975 18136 7987 18139
rect 8128 18136 8156 18176
rect 8297 18173 8309 18176
rect 8343 18173 8355 18207
rect 8297 18167 8355 18173
rect 15378 18164 15384 18216
rect 15436 18164 15442 18216
rect 15488 18204 15516 18244
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 18046 18232 18052 18284
rect 18104 18272 18110 18284
rect 18141 18275 18199 18281
rect 18141 18272 18153 18275
rect 18104 18244 18153 18272
rect 18104 18232 18110 18244
rect 18141 18241 18153 18244
rect 18187 18272 18199 18275
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 18187 18244 18245 18272
rect 18187 18241 18199 18244
rect 18141 18235 18199 18241
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 15565 18207 15623 18213
rect 15488 18176 15525 18204
rect 7975 18108 8156 18136
rect 15497 18136 15525 18176
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 15654 18204 15660 18216
rect 15611 18176 15660 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 15654 18164 15660 18176
rect 15712 18164 15718 18216
rect 15497 18108 15608 18136
rect 7975 18105 7987 18108
rect 7929 18099 7987 18105
rect 9766 18068 9772 18080
rect 7576 18040 9772 18068
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 14001 18071 14059 18077
rect 14001 18037 14013 18071
rect 14047 18068 14059 18071
rect 14090 18068 14096 18080
rect 14047 18040 14096 18068
rect 14047 18037 14059 18040
rect 14001 18031 14059 18037
rect 14090 18028 14096 18040
rect 14148 18068 14154 18080
rect 14642 18068 14648 18080
rect 14148 18040 14648 18068
rect 14148 18028 14154 18040
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 15580 18077 15608 18108
rect 16316 18108 16988 18136
rect 16316 18077 16344 18108
rect 16960 18080 16988 18108
rect 15565 18071 15623 18077
rect 15565 18037 15577 18071
rect 15611 18037 15623 18071
rect 15565 18031 15623 18037
rect 16301 18071 16359 18077
rect 16301 18037 16313 18071
rect 16347 18037 16359 18071
rect 16301 18031 16359 18037
rect 16485 18071 16543 18077
rect 16485 18037 16497 18071
rect 16531 18068 16543 18071
rect 16666 18068 16672 18080
rect 16531 18040 16672 18068
rect 16531 18037 16543 18040
rect 16485 18031 16543 18037
rect 16666 18028 16672 18040
rect 16724 18028 16730 18080
rect 16942 18028 16948 18080
rect 17000 18028 17006 18080
rect 1104 17978 20792 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 10214 17978
rect 10266 17926 10278 17978
rect 10330 17926 10342 17978
rect 10394 17926 10406 17978
rect 10458 17926 10470 17978
rect 10522 17926 16214 17978
rect 16266 17926 16278 17978
rect 16330 17926 16342 17978
rect 16394 17926 16406 17978
rect 16458 17926 16470 17978
rect 16522 17926 20792 17978
rect 1104 17904 20792 17926
rect 9306 17824 9312 17876
rect 9364 17864 9370 17876
rect 9677 17867 9735 17873
rect 9677 17864 9689 17867
rect 9364 17836 9689 17864
rect 9364 17824 9370 17836
rect 9677 17833 9689 17836
rect 9723 17833 9735 17867
rect 9677 17827 9735 17833
rect 9401 17799 9459 17805
rect 9401 17765 9413 17799
rect 9447 17765 9459 17799
rect 9401 17759 9459 17765
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17728 1731 17731
rect 1854 17728 1860 17740
rect 1719 17700 1860 17728
rect 1719 17697 1731 17700
rect 1673 17691 1731 17697
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2130 17728 2136 17740
rect 1995 17700 2136 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 2130 17688 2136 17700
rect 2188 17688 2194 17740
rect 4157 17731 4215 17737
rect 4157 17697 4169 17731
rect 4203 17728 4215 17731
rect 4706 17728 4712 17740
rect 4203 17700 4712 17728
rect 4203 17697 4215 17700
rect 4157 17691 4215 17697
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 5629 17731 5687 17737
rect 4856 17700 5580 17728
rect 4856 17688 4862 17700
rect 1578 17620 1584 17672
rect 1636 17620 1642 17672
rect 3881 17663 3939 17669
rect 3881 17629 3893 17663
rect 3927 17629 3939 17663
rect 3881 17623 3939 17629
rect 3896 17592 3924 17623
rect 3896 17564 4200 17592
rect 2958 17484 2964 17536
rect 3016 17524 3022 17536
rect 3237 17527 3295 17533
rect 3237 17524 3249 17527
rect 3016 17496 3249 17524
rect 3016 17484 3022 17496
rect 3237 17493 3249 17496
rect 3283 17524 3295 17527
rect 4062 17524 4068 17536
rect 3283 17496 4068 17524
rect 3283 17493 3295 17496
rect 3237 17487 3295 17493
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 4172 17524 4200 17564
rect 4798 17552 4804 17604
rect 4856 17552 4862 17604
rect 5552 17592 5580 17700
rect 5629 17697 5641 17731
rect 5675 17728 5687 17731
rect 6089 17731 6147 17737
rect 6089 17728 6101 17731
rect 5675 17700 6101 17728
rect 5675 17697 5687 17700
rect 5629 17691 5687 17697
rect 6089 17697 6101 17700
rect 6135 17697 6147 17731
rect 9416 17728 9444 17759
rect 6089 17691 6147 17697
rect 8772 17700 9444 17728
rect 9692 17728 9720 17827
rect 13722 17824 13728 17876
rect 13780 17864 13786 17876
rect 13817 17867 13875 17873
rect 13817 17864 13829 17867
rect 13780 17836 13829 17864
rect 13780 17824 13786 17836
rect 13817 17833 13829 17836
rect 13863 17833 13875 17867
rect 13817 17827 13875 17833
rect 14182 17824 14188 17876
rect 14240 17824 14246 17876
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 15841 17867 15899 17873
rect 15436 17836 15608 17864
rect 15436 17824 15442 17836
rect 15580 17737 15608 17836
rect 15841 17833 15853 17867
rect 15887 17864 15899 17867
rect 16114 17864 16120 17876
rect 15887 17836 16120 17864
rect 15887 17833 15899 17836
rect 15841 17827 15899 17833
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18049 17867 18107 17873
rect 18049 17864 18061 17867
rect 18012 17836 18061 17864
rect 18012 17824 18018 17836
rect 18049 17833 18061 17836
rect 18095 17833 18107 17867
rect 18049 17827 18107 17833
rect 15565 17731 15623 17737
rect 9692 17700 10180 17728
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 8772 17669 8800 17700
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17629 8631 17663
rect 8573 17623 8631 17629
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17629 8815 17663
rect 8757 17623 8815 17629
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17660 9183 17663
rect 9306 17660 9312 17672
rect 9171 17632 9312 17660
rect 9171 17629 9183 17632
rect 9125 17623 9183 17629
rect 6546 17592 6552 17604
rect 5552 17564 6552 17592
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 8588 17592 8616 17623
rect 9306 17620 9312 17632
rect 9364 17620 9370 17672
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17660 9459 17663
rect 9447 17632 10088 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 9692 17601 9720 17632
rect 9661 17595 9720 17601
rect 8588 17564 9536 17592
rect 9508 17536 9536 17564
rect 9661 17561 9673 17595
rect 9707 17564 9720 17595
rect 9707 17561 9719 17564
rect 9661 17555 9719 17561
rect 9766 17552 9772 17604
rect 9824 17592 9830 17604
rect 9861 17595 9919 17601
rect 9861 17592 9873 17595
rect 9824 17564 9873 17592
rect 9824 17552 9830 17564
rect 9861 17561 9873 17564
rect 9907 17592 9919 17595
rect 9953 17595 10011 17601
rect 9953 17592 9965 17595
rect 9907 17564 9965 17592
rect 9907 17561 9919 17564
rect 9861 17555 9919 17561
rect 9953 17561 9965 17564
rect 9999 17561 10011 17595
rect 9953 17555 10011 17561
rect 5810 17524 5816 17536
rect 4172 17496 5816 17524
rect 5810 17484 5816 17496
rect 5868 17484 5874 17536
rect 7558 17484 7564 17536
rect 7616 17484 7622 17536
rect 8662 17484 8668 17536
rect 8720 17484 8726 17536
rect 9217 17527 9275 17533
rect 9217 17493 9229 17527
rect 9263 17524 9275 17527
rect 9398 17524 9404 17536
rect 9263 17496 9404 17524
rect 9263 17493 9275 17496
rect 9217 17487 9275 17493
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 9490 17484 9496 17536
rect 9548 17484 9554 17536
rect 10060 17524 10088 17632
rect 10152 17601 10180 17700
rect 15565 17697 15577 17731
rect 15611 17697 15623 17731
rect 15565 17691 15623 17697
rect 18046 17688 18052 17740
rect 18104 17728 18110 17740
rect 18509 17731 18567 17737
rect 18509 17728 18521 17731
rect 18104 17700 18521 17728
rect 18104 17688 18110 17700
rect 18509 17697 18521 17700
rect 18555 17697 18567 17731
rect 19794 17728 19800 17740
rect 18509 17691 18567 17697
rect 19536 17700 19800 17728
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10367 17632 11100 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 10137 17595 10195 17601
rect 10137 17561 10149 17595
rect 10183 17561 10195 17595
rect 10137 17555 10195 17561
rect 10229 17595 10287 17601
rect 10229 17561 10241 17595
rect 10275 17592 10287 17595
rect 10275 17564 10364 17592
rect 10275 17561 10287 17564
rect 10229 17555 10287 17561
rect 10336 17536 10364 17564
rect 11072 17536 11100 17632
rect 14366 17620 14372 17672
rect 14424 17660 14430 17672
rect 15298 17663 15356 17669
rect 15298 17660 15310 17663
rect 14424 17632 15310 17660
rect 14424 17620 14430 17632
rect 15298 17629 15310 17632
rect 15344 17660 15356 17663
rect 15654 17660 15660 17672
rect 15344 17632 15660 17660
rect 15344 17629 15356 17632
rect 15298 17623 15356 17629
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 16942 17620 16948 17672
rect 17000 17669 17006 17672
rect 19536 17669 19564 17700
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 17000 17660 17012 17669
rect 17221 17663 17279 17669
rect 17000 17632 17045 17660
rect 17000 17623 17012 17632
rect 17221 17629 17233 17663
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 17000 17620 17006 17623
rect 16666 17552 16672 17604
rect 16724 17552 16730 17604
rect 16850 17552 16856 17604
rect 16908 17592 16914 17604
rect 17236 17592 17264 17623
rect 19610 17620 19616 17672
rect 19668 17620 19674 17672
rect 19702 17620 19708 17672
rect 19760 17620 19766 17672
rect 16908 17564 17264 17592
rect 17865 17595 17923 17601
rect 16908 17552 16914 17564
rect 17865 17561 17877 17595
rect 17911 17561 17923 17595
rect 17865 17555 17923 17561
rect 18081 17595 18139 17601
rect 18081 17561 18093 17595
rect 18127 17592 18139 17595
rect 19245 17595 19303 17601
rect 19245 17592 19257 17595
rect 18127 17564 19257 17592
rect 18127 17561 18139 17564
rect 18081 17555 18139 17561
rect 19245 17561 19257 17564
rect 19291 17561 19303 17595
rect 19245 17555 19303 17561
rect 19429 17595 19487 17601
rect 19429 17561 19441 17595
rect 19475 17592 19487 17595
rect 19720 17592 19748 17620
rect 19475 17564 19748 17592
rect 19475 17561 19487 17564
rect 19429 17555 19487 17561
rect 10318 17524 10324 17536
rect 10060 17496 10324 17524
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 10502 17484 10508 17536
rect 10560 17484 10566 17536
rect 11054 17484 11060 17536
rect 11112 17484 11118 17536
rect 16684 17524 16712 17552
rect 17880 17524 17908 17555
rect 19794 17552 19800 17604
rect 19852 17552 19858 17604
rect 16684 17496 17908 17524
rect 18230 17484 18236 17536
rect 18288 17484 18294 17536
rect 1104 17434 20792 17456
rect 1104 17382 7214 17434
rect 7266 17382 7278 17434
rect 7330 17382 7342 17434
rect 7394 17382 7406 17434
rect 7458 17382 7470 17434
rect 7522 17382 13214 17434
rect 13266 17382 13278 17434
rect 13330 17382 13342 17434
rect 13394 17382 13406 17434
rect 13458 17382 13470 17434
rect 13522 17382 19214 17434
rect 19266 17382 19278 17434
rect 19330 17382 19342 17434
rect 19394 17382 19406 17434
rect 19458 17382 19470 17434
rect 19522 17382 20792 17434
rect 1104 17360 20792 17382
rect 5166 17280 5172 17332
rect 5224 17280 5230 17332
rect 6546 17280 6552 17332
rect 6604 17280 6610 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 8720 17292 9076 17320
rect 8720 17280 8726 17292
rect 3504 17255 3562 17261
rect 1688 17224 2774 17252
rect 1688 17193 1716 17224
rect 1946 17193 1952 17196
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 1940 17147 1952 17193
rect 1946 17144 1952 17147
rect 2004 17144 2010 17196
rect 2746 17116 2774 17224
rect 3504 17221 3516 17255
rect 3550 17252 3562 17255
rect 3602 17252 3608 17264
rect 3550 17224 3608 17252
rect 3550 17221 3562 17224
rect 3504 17215 3562 17221
rect 3602 17212 3608 17224
rect 3660 17212 3666 17264
rect 6564 17252 6592 17280
rect 9048 17261 9076 17292
rect 10318 17280 10324 17332
rect 10376 17320 10382 17332
rect 10505 17323 10563 17329
rect 10505 17320 10517 17323
rect 10376 17292 10517 17320
rect 10376 17280 10382 17292
rect 10505 17289 10517 17292
rect 10551 17289 10563 17323
rect 10505 17283 10563 17289
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 12492 17292 12541 17320
rect 12492 17280 12498 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 12529 17283 12587 17289
rect 15378 17280 15384 17332
rect 15436 17320 15442 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 15436 17292 15577 17320
rect 15436 17280 15442 17292
rect 15565 17289 15577 17292
rect 15611 17320 15623 17323
rect 16850 17320 16856 17332
rect 15611 17292 16856 17320
rect 15611 17289 15623 17292
rect 15565 17283 15623 17289
rect 16850 17280 16856 17292
rect 16908 17320 16914 17332
rect 18046 17320 18052 17332
rect 16908 17292 18052 17320
rect 16908 17280 16914 17292
rect 18046 17280 18052 17292
rect 18104 17320 18110 17332
rect 18104 17292 19748 17320
rect 18104 17280 18110 17292
rect 9033 17255 9091 17261
rect 5000 17224 5672 17252
rect 6564 17224 7590 17252
rect 5000 17196 5028 17224
rect 4982 17144 4988 17196
rect 5040 17144 5046 17196
rect 5166 17144 5172 17196
rect 5224 17184 5230 17196
rect 5644 17193 5672 17224
rect 9033 17221 9045 17255
rect 9079 17221 9091 17255
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 9033 17215 9091 17221
rect 10796 17224 10977 17252
rect 5353 17187 5411 17193
rect 5353 17184 5365 17187
rect 5224 17156 5365 17184
rect 5224 17144 5230 17156
rect 5353 17153 5365 17156
rect 5399 17153 5411 17187
rect 5353 17147 5411 17153
rect 5537 17187 5595 17193
rect 5537 17153 5549 17187
rect 5583 17153 5595 17187
rect 5537 17147 5595 17153
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 2958 17116 2964 17128
rect 2746 17088 2964 17116
rect 2958 17076 2964 17088
rect 3016 17116 3022 17128
rect 3237 17119 3295 17125
rect 3237 17116 3249 17119
rect 3016 17088 3249 17116
rect 3016 17076 3022 17088
rect 3237 17085 3249 17088
rect 3283 17085 3295 17119
rect 3237 17079 3295 17085
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17085 4859 17119
rect 5552 17116 5580 17147
rect 5810 17144 5816 17196
rect 5868 17184 5874 17196
rect 5868 17156 6868 17184
rect 5868 17144 5874 17156
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 5552 17088 5733 17116
rect 4801 17079 4859 17085
rect 5721 17085 5733 17088
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 3050 16940 3056 16992
rect 3108 16940 3114 16992
rect 3252 16980 3280 17079
rect 4816 17048 4844 17079
rect 5828 17048 5856 17144
rect 6840 17125 6868 17156
rect 10042 17144 10048 17196
rect 10100 17184 10106 17196
rect 10100 17156 10166 17184
rect 10100 17144 10106 17156
rect 10502 17144 10508 17196
rect 10560 17184 10566 17196
rect 10796 17193 10824 17224
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 10965 17215 11023 17221
rect 13722 17212 13728 17264
rect 13780 17212 13786 17264
rect 13940 17255 13998 17261
rect 13940 17221 13952 17255
rect 13986 17252 13998 17255
rect 14090 17252 14096 17264
rect 13986 17224 14096 17252
rect 13986 17221 13998 17224
rect 13940 17215 13998 17221
rect 14090 17212 14096 17224
rect 14148 17212 14154 17264
rect 19460 17255 19518 17261
rect 19460 17221 19472 17255
rect 19506 17252 19518 17255
rect 19610 17252 19616 17264
rect 19506 17224 19616 17252
rect 19506 17221 19518 17224
rect 19460 17215 19518 17221
rect 19610 17212 19616 17224
rect 19668 17212 19674 17264
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10560 17156 10609 17184
rect 10560 17144 10566 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17153 10931 17187
rect 10873 17147 10931 17153
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17116 7159 17119
rect 7558 17116 7564 17128
rect 7147 17088 7564 17116
rect 7147 17085 7159 17088
rect 7101 17079 7159 17085
rect 4816 17020 5856 17048
rect 3510 16980 3516 16992
rect 3252 16952 3516 16980
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 4614 16940 4620 16992
rect 4672 16940 4678 16992
rect 5534 16940 5540 16992
rect 5592 16940 5598 16992
rect 6840 16980 6868 17079
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 8570 17076 8576 17128
rect 8628 17116 8634 17128
rect 8757 17119 8815 17125
rect 8757 17116 8769 17119
rect 8628 17088 8769 17116
rect 8628 17076 8634 17088
rect 8757 17085 8769 17088
rect 8803 17085 8815 17119
rect 8757 17079 8815 17085
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 10888 17116 10916 17147
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 12342 17184 12348 17196
rect 11112 17156 12348 17184
rect 11112 17144 11118 17156
rect 12342 17144 12348 17156
rect 12400 17144 12406 17196
rect 13740 17184 13768 17212
rect 19720 17193 19748 17292
rect 14185 17187 14243 17193
rect 14185 17184 14197 17187
rect 13740 17156 14197 17184
rect 14185 17153 14197 17156
rect 14231 17153 14243 17187
rect 14185 17147 14243 17153
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 9548 17088 10916 17116
rect 9548 17076 9554 17088
rect 7098 16980 7104 16992
rect 6840 16952 7104 16980
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 8573 16983 8631 16989
rect 8573 16949 8585 16983
rect 8619 16980 8631 16983
rect 8662 16980 8668 16992
rect 8619 16952 8668 16980
rect 8619 16949 8631 16952
rect 8573 16943 8631 16949
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 10781 16983 10839 16989
rect 10781 16949 10793 16983
rect 10827 16980 10839 16983
rect 10870 16980 10876 16992
rect 10827 16952 10876 16980
rect 10827 16949 10839 16952
rect 10781 16943 10839 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 12802 16940 12808 16992
rect 12860 16940 12866 16992
rect 18322 16940 18328 16992
rect 18380 16980 18386 16992
rect 19794 16980 19800 16992
rect 18380 16952 19800 16980
rect 18380 16940 18386 16952
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 1104 16890 20792 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 10214 16890
rect 10266 16838 10278 16890
rect 10330 16838 10342 16890
rect 10394 16838 10406 16890
rect 10458 16838 10470 16890
rect 10522 16838 16214 16890
rect 16266 16838 16278 16890
rect 16330 16838 16342 16890
rect 16394 16838 16406 16890
rect 16458 16838 16470 16890
rect 16522 16838 20792 16890
rect 1104 16816 20792 16838
rect 3510 16776 3516 16788
rect 1872 16748 3516 16776
rect 1670 16600 1676 16652
rect 1728 16600 1734 16652
rect 1872 16649 1900 16748
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 3602 16736 3608 16788
rect 3660 16736 3666 16788
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 3973 16779 4031 16785
rect 3973 16776 3985 16779
rect 3936 16748 3985 16776
rect 3936 16736 3942 16748
rect 3973 16745 3985 16748
rect 4019 16745 4031 16779
rect 3973 16739 4031 16745
rect 4157 16779 4215 16785
rect 4157 16745 4169 16779
rect 4203 16776 4215 16779
rect 4982 16776 4988 16788
rect 4203 16748 4988 16776
rect 4203 16745 4215 16748
rect 4157 16739 4215 16745
rect 3421 16711 3479 16717
rect 3421 16677 3433 16711
rect 3467 16708 3479 16711
rect 3620 16708 3648 16736
rect 4172 16708 4200 16739
rect 4982 16736 4988 16748
rect 5040 16736 5046 16788
rect 10870 16785 10876 16788
rect 5629 16779 5687 16785
rect 5629 16745 5641 16779
rect 5675 16776 5687 16779
rect 10854 16779 10876 16785
rect 5675 16748 8616 16776
rect 5675 16745 5687 16748
rect 5629 16739 5687 16745
rect 3467 16680 3648 16708
rect 3804 16680 4200 16708
rect 4525 16711 4583 16717
rect 3467 16677 3479 16680
rect 3421 16671 3479 16677
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16609 1915 16643
rect 3694 16640 3700 16652
rect 1857 16603 1915 16609
rect 3436 16612 3700 16640
rect 2130 16581 2136 16584
rect 2124 16572 2136 16581
rect 2091 16544 2136 16572
rect 2124 16535 2136 16544
rect 2130 16532 2136 16535
rect 2188 16532 2194 16584
rect 3436 16581 3464 16612
rect 3694 16600 3700 16612
rect 3752 16600 3758 16652
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 3804 16572 3832 16680
rect 4525 16677 4537 16711
rect 4571 16677 4583 16711
rect 4525 16671 4583 16677
rect 3970 16600 3976 16652
rect 4028 16640 4034 16652
rect 4540 16640 4568 16671
rect 5736 16649 5764 16748
rect 8588 16652 8616 16748
rect 10854 16745 10866 16779
rect 10854 16739 10876 16745
rect 10870 16736 10876 16739
rect 10928 16736 10934 16788
rect 12342 16736 12348 16788
rect 12400 16736 12406 16788
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 13780 16748 14381 16776
rect 13780 16736 13786 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 14369 16739 14427 16745
rect 4028 16612 4568 16640
rect 5721 16643 5779 16649
rect 4028 16600 4034 16612
rect 5721 16609 5733 16643
rect 5767 16609 5779 16643
rect 5721 16603 5779 16609
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 8665 16643 8723 16649
rect 8665 16640 8677 16643
rect 8628 16612 8677 16640
rect 8628 16600 8634 16612
rect 8665 16609 8677 16612
rect 8711 16640 8723 16643
rect 10505 16643 10563 16649
rect 10505 16640 10517 16643
rect 8711 16612 10517 16640
rect 8711 16609 8723 16612
rect 8665 16603 8723 16609
rect 10505 16609 10517 16612
rect 10551 16640 10563 16643
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 10551 16612 10609 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 10597 16609 10609 16612
rect 10643 16640 10655 16643
rect 10962 16640 10968 16652
rect 10643 16612 10968 16640
rect 10643 16609 10655 16612
rect 10597 16603 10655 16609
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 14384 16640 14412 16739
rect 15194 16736 15200 16788
rect 15252 16736 15258 16788
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 17405 16779 17463 16785
rect 17405 16776 17417 16779
rect 16908 16748 17417 16776
rect 16908 16736 16914 16748
rect 17405 16745 17417 16748
rect 17451 16745 17463 16779
rect 17405 16739 17463 16745
rect 15212 16708 15240 16736
rect 15212 16680 15608 16708
rect 15580 16649 15608 16680
rect 15105 16643 15163 16649
rect 14384 16612 15056 16640
rect 15028 16584 15056 16612
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15381 16643 15439 16649
rect 15381 16640 15393 16643
rect 15151 16612 15393 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 15381 16609 15393 16612
rect 15427 16609 15439 16643
rect 15381 16603 15439 16609
rect 15565 16643 15623 16649
rect 15565 16609 15577 16643
rect 15611 16609 15623 16643
rect 15565 16603 15623 16609
rect 15841 16643 15899 16649
rect 15841 16609 15853 16643
rect 15887 16640 15899 16643
rect 17126 16640 17132 16652
rect 15887 16612 17132 16640
rect 15887 16609 15899 16612
rect 15841 16603 15899 16609
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 17420 16640 17448 16739
rect 17589 16643 17647 16649
rect 17589 16640 17601 16643
rect 17420 16612 17601 16640
rect 17589 16609 17601 16612
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 3651 16544 3832 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 3878 16532 3884 16584
rect 3936 16572 3942 16584
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 3936 16544 4261 16572
rect 3936 16532 3942 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 5977 16575 6035 16581
rect 5977 16572 5989 16575
rect 5592 16544 5989 16572
rect 5592 16532 5598 16544
rect 5977 16541 5989 16544
rect 6023 16541 6035 16575
rect 5977 16535 6035 16541
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14424 16544 14565 16572
rect 14424 16532 14430 16544
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 15197 16575 15255 16581
rect 15197 16541 15209 16575
rect 15243 16572 15255 16575
rect 15470 16572 15476 16584
rect 15243 16544 15476 16572
rect 15243 16541 15255 16544
rect 15197 16535 15255 16541
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 15654 16532 15660 16584
rect 15712 16532 15718 16584
rect 17856 16575 17914 16581
rect 17856 16541 17868 16575
rect 17902 16572 17914 16575
rect 18322 16572 18328 16584
rect 17902 16544 18328 16572
rect 17902 16541 17914 16544
rect 17856 16535 17914 16541
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 20254 16532 20260 16584
rect 20312 16532 20318 16584
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 1489 16507 1547 16513
rect 1489 16504 1501 16507
rect 992 16476 1501 16504
rect 992 16464 998 16476
rect 1489 16473 1501 16476
rect 1535 16473 1547 16507
rect 1489 16467 1547 16473
rect 1578 16464 1584 16516
rect 1636 16504 1642 16516
rect 3050 16504 3056 16516
rect 1636 16476 3056 16504
rect 1636 16464 1642 16476
rect 3050 16464 3056 16476
rect 3108 16504 3114 16516
rect 3789 16507 3847 16513
rect 3789 16504 3801 16507
rect 3108 16476 3801 16504
rect 3108 16464 3114 16476
rect 3789 16473 3801 16476
rect 3835 16504 3847 16507
rect 4341 16507 4399 16513
rect 4341 16504 4353 16507
rect 3835 16476 4353 16504
rect 3835 16473 3847 16476
rect 3789 16467 3847 16473
rect 4341 16473 4353 16476
rect 4387 16473 4399 16507
rect 4341 16467 4399 16473
rect 4525 16507 4583 16513
rect 4525 16473 4537 16507
rect 4571 16504 4583 16507
rect 4614 16504 4620 16516
rect 4571 16476 4620 16504
rect 4571 16473 4583 16476
rect 4525 16467 4583 16473
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 3326 16436 3332 16448
rect 3283 16408 3332 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 3326 16396 3332 16408
rect 3384 16436 3390 16448
rect 3878 16436 3884 16448
rect 3384 16408 3884 16436
rect 3384 16396 3390 16408
rect 3878 16396 3884 16408
rect 3936 16396 3942 16448
rect 3970 16396 3976 16448
rect 4028 16445 4034 16448
rect 4028 16439 4047 16445
rect 4035 16436 4047 16439
rect 4540 16436 4568 16467
rect 4614 16464 4620 16476
rect 4672 16464 4678 16516
rect 14921 16507 14979 16513
rect 14921 16504 14933 16507
rect 12098 16476 12434 16504
rect 4035 16408 4568 16436
rect 4035 16405 4047 16408
rect 4028 16399 4047 16405
rect 4028 16396 4034 16399
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 7834 16436 7840 16448
rect 7156 16408 7840 16436
rect 7156 16396 7162 16408
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 12406 16436 12434 16476
rect 14660 16476 14933 16504
rect 13078 16436 13084 16448
rect 12406 16408 13084 16436
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 14458 16396 14464 16448
rect 14516 16436 14522 16448
rect 14660 16436 14688 16476
rect 14921 16473 14933 16476
rect 14967 16473 14979 16507
rect 14921 16467 14979 16473
rect 15286 16464 15292 16516
rect 15344 16464 15350 16516
rect 15488 16504 15516 16532
rect 16022 16504 16028 16516
rect 15488 16476 16028 16504
rect 16022 16464 16028 16476
rect 16080 16464 16086 16516
rect 20272 16504 20300 16532
rect 17880 16476 20300 16504
rect 17880 16448 17908 16476
rect 14516 16408 14688 16436
rect 14516 16396 14522 16408
rect 14734 16396 14740 16448
rect 14792 16396 14798 16448
rect 14826 16396 14832 16448
rect 14884 16396 14890 16448
rect 17862 16396 17868 16448
rect 17920 16396 17926 16448
rect 18966 16396 18972 16448
rect 19024 16396 19030 16448
rect 1104 16346 20792 16368
rect 1104 16294 7214 16346
rect 7266 16294 7278 16346
rect 7330 16294 7342 16346
rect 7394 16294 7406 16346
rect 7458 16294 7470 16346
rect 7522 16294 13214 16346
rect 13266 16294 13278 16346
rect 13330 16294 13342 16346
rect 13394 16294 13406 16346
rect 13458 16294 13470 16346
rect 13522 16294 19214 16346
rect 19266 16294 19278 16346
rect 19330 16294 19342 16346
rect 19394 16294 19406 16346
rect 19458 16294 19470 16346
rect 19522 16294 20792 16346
rect 1104 16272 20792 16294
rect 1946 16192 1952 16244
rect 2004 16192 2010 16244
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12713 16235 12771 16241
rect 12713 16232 12725 16235
rect 12492 16204 12725 16232
rect 12492 16192 12498 16204
rect 12713 16201 12725 16204
rect 12759 16201 12771 16235
rect 12713 16195 12771 16201
rect 14277 16235 14335 16241
rect 14277 16201 14289 16235
rect 14323 16232 14335 16235
rect 14826 16232 14832 16244
rect 14323 16204 14832 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 1578 16124 1584 16176
rect 1636 16124 1642 16176
rect 10594 16164 10600 16176
rect 10520 16136 10600 16164
rect 1596 16096 1624 16124
rect 2038 16096 2044 16108
rect 1596 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10520 16105 10548 16136
rect 10594 16124 10600 16136
rect 10652 16124 10658 16176
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10192 16068 10333 16096
rect 10192 16056 10198 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 10505 16099 10563 16105
rect 10505 16065 10517 16099
rect 10551 16065 10563 16099
rect 12728 16096 12756 16195
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 15286 16192 15292 16244
rect 15344 16232 15350 16244
rect 15930 16232 15936 16244
rect 15344 16204 15936 16232
rect 15344 16192 15350 16204
rect 15930 16192 15936 16204
rect 15988 16232 15994 16244
rect 16393 16235 16451 16241
rect 16393 16232 16405 16235
rect 15988 16204 16405 16232
rect 15988 16192 15994 16204
rect 16393 16201 16405 16204
rect 16439 16201 16451 16235
rect 16393 16195 16451 16201
rect 17236 16204 18460 16232
rect 12802 16124 12808 16176
rect 12860 16164 12866 16176
rect 13142 16167 13200 16173
rect 13142 16164 13154 16167
rect 12860 16136 13154 16164
rect 12860 16124 12866 16136
rect 13142 16133 13154 16136
rect 13188 16164 13200 16167
rect 14458 16164 14464 16176
rect 13188 16136 14464 16164
rect 13188 16133 13200 16136
rect 13142 16127 13200 16133
rect 14458 16124 14464 16136
rect 14516 16124 14522 16176
rect 14844 16164 14872 16192
rect 14660 16136 14872 16164
rect 12897 16099 12955 16105
rect 12897 16096 12909 16099
rect 12728 16068 12909 16096
rect 10505 16059 10563 16065
rect 12897 16065 12909 16068
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 14366 16056 14372 16108
rect 14424 16056 14430 16108
rect 14660 16105 14688 16136
rect 16022 16124 16028 16176
rect 16080 16164 16086 16176
rect 17236 16173 17264 16204
rect 17221 16167 17279 16173
rect 17221 16164 17233 16167
rect 16080 16136 17233 16164
rect 16080 16124 16086 16136
rect 17221 16133 17233 16136
rect 17267 16133 17279 16167
rect 17221 16127 17279 16133
rect 17589 16167 17647 16173
rect 17589 16133 17601 16167
rect 17635 16164 17647 16167
rect 18138 16164 18144 16176
rect 17635 16136 18144 16164
rect 17635 16133 17647 16136
rect 17589 16127 17647 16133
rect 18138 16124 18144 16136
rect 18196 16124 18202 16176
rect 18230 16124 18236 16176
rect 18288 16124 18294 16176
rect 18432 16173 18460 16204
rect 18417 16167 18475 16173
rect 18417 16133 18429 16167
rect 18463 16133 18475 16167
rect 18417 16127 18475 16133
rect 14645 16099 14703 16105
rect 14645 16065 14657 16099
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16096 14795 16099
rect 15269 16099 15327 16105
rect 15269 16096 15281 16099
rect 14783 16068 15281 16096
rect 14783 16065 14795 16068
rect 14737 16059 14795 16065
rect 15269 16065 15281 16068
rect 15315 16065 15327 16099
rect 15269 16059 15327 16065
rect 17957 16099 18015 16105
rect 17957 16065 17969 16099
rect 18003 16065 18015 16099
rect 17957 16059 18015 16065
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18248 16096 18276 16124
rect 18095 16068 18276 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 14384 16028 14412 16056
rect 14752 16028 14780 16059
rect 14384 16000 14780 16028
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 17972 16028 18000 16059
rect 18966 16056 18972 16108
rect 19024 16096 19030 16108
rect 20082 16099 20140 16105
rect 20082 16096 20094 16099
rect 19024 16068 20094 16096
rect 19024 16056 19030 16068
rect 20082 16065 20094 16068
rect 20128 16065 20140 16099
rect 20082 16059 20140 16065
rect 20346 16056 20352 16108
rect 20404 16056 20410 16108
rect 17604 16000 18000 16028
rect 14734 15960 14740 15972
rect 14660 15932 14740 15960
rect 3510 15852 3516 15904
rect 3568 15852 3574 15904
rect 10413 15895 10471 15901
rect 10413 15861 10425 15895
rect 10459 15892 10471 15895
rect 10594 15892 10600 15904
rect 10459 15864 10600 15892
rect 10459 15861 10471 15864
rect 10413 15855 10471 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11054 15852 11060 15904
rect 11112 15852 11118 15904
rect 14660 15901 14688 15932
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 17310 15920 17316 15972
rect 17368 15960 17374 15972
rect 17604 15969 17632 16000
rect 18230 15988 18236 16040
rect 18288 15988 18294 16040
rect 18325 16031 18383 16037
rect 18325 15997 18337 16031
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 17589 15963 17647 15969
rect 17368 15932 17540 15960
rect 17368 15920 17374 15932
rect 14645 15895 14703 15901
rect 14645 15861 14657 15895
rect 14691 15861 14703 15895
rect 14645 15855 14703 15861
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 15378 15892 15384 15904
rect 14967 15864 15384 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 17402 15852 17408 15904
rect 17460 15852 17466 15904
rect 17512 15892 17540 15932
rect 17589 15929 17601 15963
rect 17635 15929 17647 15963
rect 18340 15960 18368 15991
rect 17589 15923 17647 15929
rect 17696 15932 18368 15960
rect 17696 15892 17724 15932
rect 17512 15864 17724 15892
rect 17770 15852 17776 15904
rect 17828 15852 17834 15904
rect 18690 15852 18696 15904
rect 18748 15852 18754 15904
rect 18969 15895 19027 15901
rect 18969 15861 18981 15895
rect 19015 15892 19027 15895
rect 19610 15892 19616 15904
rect 19015 15864 19616 15892
rect 19015 15861 19027 15864
rect 18969 15855 19027 15861
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 1104 15802 20792 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 10214 15802
rect 10266 15750 10278 15802
rect 10330 15750 10342 15802
rect 10394 15750 10406 15802
rect 10458 15750 10470 15802
rect 10522 15750 16214 15802
rect 16266 15750 16278 15802
rect 16330 15750 16342 15802
rect 16394 15750 16406 15802
rect 16458 15750 16470 15802
rect 16522 15750 20792 15802
rect 1104 15728 20792 15750
rect 10594 15648 10600 15700
rect 10652 15648 10658 15700
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 11146 15688 11152 15700
rect 10744 15660 11152 15688
rect 10744 15648 10750 15660
rect 11146 15648 11152 15660
rect 11204 15688 11210 15700
rect 11790 15688 11796 15700
rect 11204 15660 11796 15688
rect 11204 15648 11210 15660
rect 11790 15648 11796 15660
rect 11848 15648 11854 15700
rect 13722 15648 13728 15700
rect 13780 15688 13786 15700
rect 13817 15691 13875 15697
rect 13817 15688 13829 15691
rect 13780 15660 13829 15688
rect 13780 15648 13786 15660
rect 13817 15657 13829 15660
rect 13863 15657 13875 15691
rect 13817 15651 13875 15657
rect 4341 15623 4399 15629
rect 4341 15589 4353 15623
rect 4387 15589 4399 15623
rect 4341 15583 4399 15589
rect 3326 15552 3332 15564
rect 1964 15524 3332 15552
rect 1964 15428 1992 15524
rect 3326 15512 3332 15524
rect 3384 15552 3390 15564
rect 4356 15552 4384 15583
rect 6362 15552 6368 15564
rect 3384 15524 4108 15552
rect 4356 15524 6368 15552
rect 3384 15512 3390 15524
rect 3789 15487 3847 15493
rect 3789 15453 3801 15487
rect 3835 15484 3847 15487
rect 3878 15484 3884 15496
rect 3835 15456 3884 15484
rect 3835 15453 3847 15456
rect 3789 15447 3847 15453
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 4080 15493 4108 15524
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 9953 15555 10011 15561
rect 9953 15552 9965 15555
rect 9692 15524 9965 15552
rect 4065 15487 4123 15493
rect 4065 15453 4077 15487
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 4433 15487 4491 15493
rect 4433 15484 4445 15487
rect 4264 15456 4445 15484
rect 1946 15376 1952 15428
rect 2004 15376 2010 15428
rect 3970 15416 3976 15428
rect 3804 15388 3976 15416
rect 3804 15360 3832 15388
rect 3970 15376 3976 15388
rect 4028 15376 4034 15428
rect 3786 15308 3792 15360
rect 3844 15348 3850 15360
rect 4264 15348 4292 15456
rect 4433 15453 4445 15456
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 4890 15444 4896 15496
rect 4948 15444 4954 15496
rect 9692 15493 9720 15524
rect 9953 15521 9965 15524
rect 9999 15521 10011 15555
rect 9953 15515 10011 15521
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15552 10563 15555
rect 10612 15552 10640 15648
rect 11514 15552 11520 15564
rect 10551 15524 10640 15552
rect 10980 15524 11520 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15484 9459 15487
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 9447 15456 9505 15484
rect 9447 15453 9459 15456
rect 9401 15447 9459 15453
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15484 9919 15487
rect 10520 15484 10548 15515
rect 9907 15456 10548 15484
rect 10597 15487 10655 15493
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 10597 15453 10609 15487
rect 10643 15484 10655 15487
rect 10980 15484 11008 15524
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 13832 15552 13860 15651
rect 14734 15648 14740 15700
rect 14792 15688 14798 15700
rect 14792 15660 15056 15688
rect 14792 15648 14798 15660
rect 15028 15620 15056 15660
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 15841 15691 15899 15697
rect 15841 15688 15853 15691
rect 15436 15660 15853 15688
rect 15436 15648 15442 15660
rect 15841 15657 15853 15660
rect 15887 15657 15899 15691
rect 15841 15651 15899 15657
rect 15930 15648 15936 15700
rect 15988 15648 15994 15700
rect 16945 15691 17003 15697
rect 16945 15657 16957 15691
rect 16991 15688 17003 15691
rect 17310 15688 17316 15700
rect 16991 15660 17316 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 17310 15648 17316 15660
rect 17368 15648 17374 15700
rect 17402 15648 17408 15700
rect 17460 15688 17466 15700
rect 18601 15691 18659 15697
rect 18601 15688 18613 15691
rect 17460 15660 18613 15688
rect 17460 15648 17466 15660
rect 18601 15657 18613 15660
rect 18647 15657 18659 15691
rect 18601 15651 18659 15657
rect 18874 15648 18880 15700
rect 18932 15648 18938 15700
rect 20438 15648 20444 15700
rect 20496 15648 20502 15700
rect 15470 15620 15476 15632
rect 15028 15592 15476 15620
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 15654 15580 15660 15632
rect 15712 15580 15718 15632
rect 18322 15580 18328 15632
rect 18380 15620 18386 15632
rect 19797 15623 19855 15629
rect 19797 15620 19809 15623
rect 18380 15592 19809 15620
rect 18380 15580 18386 15592
rect 19797 15589 19809 15592
rect 19843 15589 19855 15623
rect 19797 15583 19855 15589
rect 14090 15552 14096 15564
rect 13832 15524 14096 15552
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 16022 15512 16028 15564
rect 16080 15512 16086 15564
rect 19245 15555 19303 15561
rect 19245 15552 19257 15555
rect 18800 15524 19257 15552
rect 18800 15496 18828 15524
rect 19245 15521 19257 15524
rect 19291 15521 19303 15555
rect 19245 15515 19303 15521
rect 10643 15456 11008 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 11149 15487 11207 15493
rect 11149 15484 11161 15487
rect 11112 15456 11161 15484
rect 11112 15444 11118 15456
rect 11149 15453 11161 15456
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 14360 15487 14418 15493
rect 14360 15453 14372 15487
rect 14406 15484 14418 15487
rect 14826 15484 14832 15496
rect 14406 15456 14832 15484
rect 14406 15453 14418 15456
rect 14360 15447 14418 15453
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 15562 15444 15568 15496
rect 15620 15484 15626 15496
rect 15657 15487 15715 15493
rect 15657 15484 15669 15487
rect 15620 15456 15669 15484
rect 15620 15444 15626 15456
rect 15657 15453 15669 15456
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 18288 15456 18337 15484
rect 18288 15444 18294 15456
rect 18325 15453 18337 15456
rect 18371 15484 18383 15487
rect 18690 15484 18696 15496
rect 18371 15456 18696 15484
rect 18371 15453 18383 15456
rect 18325 15447 18383 15453
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 18782 15444 18788 15496
rect 18840 15444 18846 15496
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 4525 15419 4583 15425
rect 4525 15385 4537 15419
rect 4571 15416 4583 15419
rect 6178 15416 6184 15428
rect 4571 15388 6184 15416
rect 4571 15385 4583 15388
rect 4525 15379 4583 15385
rect 6178 15376 6184 15388
rect 6236 15376 6242 15428
rect 6638 15376 6644 15428
rect 6696 15376 6702 15428
rect 8018 15416 8024 15428
rect 7866 15388 8024 15416
rect 8018 15376 8024 15388
rect 8076 15376 8082 15428
rect 10137 15419 10195 15425
rect 10137 15385 10149 15419
rect 10183 15416 10195 15419
rect 10226 15416 10232 15428
rect 10183 15388 10232 15416
rect 10183 15385 10195 15388
rect 10137 15379 10195 15385
rect 10226 15376 10232 15388
rect 10284 15376 10290 15428
rect 10321 15419 10379 15425
rect 10321 15385 10333 15419
rect 10367 15416 10379 15419
rect 10686 15416 10692 15428
rect 10367 15388 10692 15416
rect 10367 15385 10379 15388
rect 10321 15379 10379 15385
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 11425 15419 11483 15425
rect 11425 15416 11437 15419
rect 10980 15388 11437 15416
rect 3844 15320 4292 15348
rect 3844 15308 3850 15320
rect 4706 15308 4712 15360
rect 4764 15308 4770 15360
rect 7650 15308 7656 15360
rect 7708 15348 7714 15360
rect 8113 15351 8171 15357
rect 8113 15348 8125 15351
rect 7708 15320 8125 15348
rect 7708 15308 7714 15320
rect 8113 15317 8125 15320
rect 8159 15317 8171 15351
rect 8113 15311 8171 15317
rect 9214 15308 9220 15360
rect 9272 15308 9278 15360
rect 10980 15357 11008 15388
rect 11425 15385 11437 15388
rect 11471 15385 11483 15419
rect 12710 15416 12716 15428
rect 12650 15388 12716 15416
rect 11425 15379 11483 15385
rect 12710 15376 12716 15388
rect 12768 15416 12774 15428
rect 12989 15419 13047 15425
rect 12989 15416 13001 15419
rect 12768 15388 13001 15416
rect 12768 15376 12774 15388
rect 12989 15385 13001 15388
rect 13035 15385 13047 15419
rect 12989 15379 13047 15385
rect 13078 15376 13084 15428
rect 13136 15416 13142 15428
rect 13357 15419 13415 15425
rect 13357 15416 13369 15419
rect 13136 15388 13369 15416
rect 13136 15376 13142 15388
rect 13357 15385 13369 15388
rect 13403 15416 13415 15419
rect 17862 15416 17868 15428
rect 13403 15388 17868 15416
rect 13403 15385 13415 15388
rect 13357 15379 13415 15385
rect 17862 15376 17868 15388
rect 17920 15376 17926 15428
rect 18080 15419 18138 15425
rect 18080 15385 18092 15419
rect 18126 15416 18138 15419
rect 18800 15416 18828 15444
rect 18126 15388 18828 15416
rect 18892 15416 18920 15447
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 19061 15487 19119 15493
rect 19061 15484 19073 15487
rect 19024 15456 19073 15484
rect 19024 15444 19030 15456
rect 19061 15453 19073 15456
rect 19107 15484 19119 15487
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 19107 15456 19625 15484
rect 19107 15453 19119 15456
rect 19061 15447 19119 15453
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 20254 15444 20260 15496
rect 20312 15444 20318 15496
rect 18892 15388 19564 15416
rect 18126 15385 18138 15388
rect 18080 15379 18138 15385
rect 10965 15351 11023 15357
rect 10965 15317 10977 15351
rect 11011 15317 11023 15351
rect 10965 15311 11023 15317
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 12897 15351 12955 15357
rect 12897 15348 12909 15351
rect 11756 15320 12909 15348
rect 11756 15308 11762 15320
rect 12897 15317 12909 15320
rect 12943 15317 12955 15351
rect 12897 15311 12955 15317
rect 16666 15308 16672 15360
rect 16724 15308 16730 15360
rect 18874 15308 18880 15360
rect 18932 15348 18938 15360
rect 19536 15357 19564 15388
rect 19429 15351 19487 15357
rect 19429 15348 19441 15351
rect 18932 15320 19441 15348
rect 18932 15308 18938 15320
rect 19429 15317 19441 15320
rect 19475 15317 19487 15351
rect 19429 15311 19487 15317
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 19610 15348 19616 15360
rect 19567 15320 19616 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 1104 15258 20792 15280
rect 1104 15206 7214 15258
rect 7266 15206 7278 15258
rect 7330 15206 7342 15258
rect 7394 15206 7406 15258
rect 7458 15206 7470 15258
rect 7522 15206 13214 15258
rect 13266 15206 13278 15258
rect 13330 15206 13342 15258
rect 13394 15206 13406 15258
rect 13458 15206 13470 15258
rect 13522 15206 19214 15258
rect 19266 15206 19278 15258
rect 19330 15206 19342 15258
rect 19394 15206 19406 15258
rect 19458 15206 19470 15258
rect 19522 15206 20792 15258
rect 1104 15184 20792 15206
rect 3789 15147 3847 15153
rect 1688 15116 3648 15144
rect 1688 15017 1716 15116
rect 1857 15079 1915 15085
rect 1857 15045 1869 15079
rect 1903 15076 1915 15079
rect 1903 15048 2084 15076
rect 1903 15045 1915 15048
rect 1857 15039 1915 15045
rect 1489 15011 1547 15017
rect 1489 14977 1501 15011
rect 1535 15008 1547 15011
rect 1673 15011 1731 15017
rect 1535 14980 1624 15008
rect 1535 14977 1547 14980
rect 1489 14971 1547 14977
rect 1486 14764 1492 14816
rect 1544 14764 1550 14816
rect 1596 14804 1624 14980
rect 1673 14977 1685 15011
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 1780 14940 1808 14971
rect 1946 14940 1952 14952
rect 1780 14912 1952 14940
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 2056 14949 2084 15048
rect 2314 15036 2320 15088
rect 2372 15036 2378 15088
rect 3620 15008 3648 15116
rect 3789 15113 3801 15147
rect 3835 15144 3847 15147
rect 4341 15147 4399 15153
rect 3835 15116 3924 15144
rect 3835 15113 3847 15116
rect 3789 15107 3847 15113
rect 3896 15085 3924 15116
rect 4341 15113 4353 15147
rect 4387 15144 4399 15147
rect 4890 15144 4896 15156
rect 4387 15116 4896 15144
rect 4387 15113 4399 15116
rect 4341 15107 4399 15113
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 6638 15104 6644 15156
rect 6696 15104 6702 15156
rect 7650 15144 7656 15156
rect 7024 15116 7656 15144
rect 3881 15079 3939 15085
rect 3881 15045 3893 15079
rect 3927 15076 3939 15079
rect 4154 15076 4160 15088
rect 3927 15048 4160 15076
rect 3927 15045 3939 15048
rect 3881 15039 3939 15045
rect 4154 15036 4160 15048
rect 4212 15036 4218 15088
rect 5258 15036 5264 15088
rect 5316 15036 5322 15088
rect 7024 15085 7052 15116
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 9214 15104 9220 15156
rect 9272 15104 9278 15156
rect 10962 15104 10968 15156
rect 11020 15144 11026 15156
rect 12069 15147 12127 15153
rect 12069 15144 12081 15147
rect 11020 15116 12081 15144
rect 11020 15104 11026 15116
rect 12069 15113 12081 15116
rect 12115 15144 12127 15147
rect 12115 15116 12434 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 7009 15079 7067 15085
rect 7009 15045 7021 15079
rect 7055 15045 7067 15079
rect 7009 15039 7067 15045
rect 8849 15079 8907 15085
rect 8849 15045 8861 15079
rect 8895 15076 8907 15079
rect 9232 15076 9260 15104
rect 11793 15079 11851 15085
rect 11793 15076 11805 15079
rect 8895 15048 9260 15076
rect 10888 15048 11805 15076
rect 8895 15045 8907 15048
rect 8849 15039 8907 15045
rect 3450 14980 3556 15008
rect 3620 14980 3924 15008
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14909 2099 14943
rect 3528 14940 3556 14980
rect 3896 14952 3924 14980
rect 6454 14968 6460 15020
rect 6512 14968 6518 15020
rect 8018 14968 8024 15020
rect 8076 15008 8082 15020
rect 8478 15008 8484 15020
rect 8076 14980 8484 15008
rect 8076 14968 8082 14980
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 8570 14968 8576 15020
rect 8628 14968 8634 15020
rect 10134 15008 10140 15020
rect 9982 14980 10140 15008
rect 10134 14968 10140 14980
rect 10192 14968 10198 15020
rect 10888 15017 10916 15048
rect 11793 15045 11805 15048
rect 11839 15076 11851 15079
rect 11839 15048 12020 15076
rect 11839 15045 11851 15048
rect 11793 15039 11851 15045
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 11057 15011 11115 15017
rect 11057 14977 11069 15011
rect 11103 15008 11115 15011
rect 11698 15008 11704 15020
rect 11103 14980 11704 15008
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 11885 15011 11943 15017
rect 11885 15008 11897 15011
rect 11808 14980 11897 15008
rect 11808 14952 11836 14980
rect 11885 14977 11897 14980
rect 11931 14977 11943 15011
rect 11885 14971 11943 14977
rect 3694 14940 3700 14952
rect 3528 14912 3700 14940
rect 2041 14903 2099 14909
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 3878 14900 3884 14952
rect 3936 14940 3942 14952
rect 4433 14943 4491 14949
rect 4433 14940 4445 14943
rect 3936 14912 4445 14940
rect 3936 14900 3942 14912
rect 4433 14909 4445 14912
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 5902 14900 5908 14952
rect 5960 14900 5966 14952
rect 6178 14900 6184 14952
rect 6236 14900 6242 14952
rect 6730 14900 6736 14952
rect 6788 14900 6794 14952
rect 10226 14900 10232 14952
rect 10284 14940 10290 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 10284 14912 10333 14940
rect 10284 14900 10290 14912
rect 10321 14909 10333 14912
rect 10367 14940 10379 14943
rect 10965 14943 11023 14949
rect 10965 14940 10977 14943
rect 10367 14912 10977 14940
rect 10367 14909 10379 14912
rect 10321 14903 10379 14909
rect 10965 14909 10977 14912
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 4157 14875 4215 14881
rect 4157 14841 4169 14875
rect 4203 14841 4215 14875
rect 4157 14835 4215 14841
rect 2130 14804 2136 14816
rect 1596 14776 2136 14804
rect 2130 14764 2136 14776
rect 2188 14804 2194 14816
rect 4172 14804 4200 14835
rect 2188 14776 4200 14804
rect 2188 14764 2194 14776
rect 7742 14764 7748 14816
rect 7800 14804 7806 14816
rect 8481 14807 8539 14813
rect 8481 14804 8493 14807
rect 7800 14776 8493 14804
rect 7800 14764 7806 14776
rect 8481 14773 8493 14776
rect 8527 14773 8539 14807
rect 10980 14804 11008 14903
rect 11146 14900 11152 14952
rect 11204 14940 11210 14952
rect 11333 14943 11391 14949
rect 11204 14912 11248 14940
rect 11204 14900 11210 14912
rect 11333 14909 11345 14943
rect 11379 14940 11391 14943
rect 11379 14912 11652 14940
rect 11379 14909 11391 14912
rect 11333 14903 11391 14909
rect 11517 14875 11575 14881
rect 11517 14841 11529 14875
rect 11563 14841 11575 14875
rect 11624 14872 11652 14912
rect 11790 14900 11796 14952
rect 11848 14900 11854 14952
rect 11992 14940 12020 15048
rect 12406 15008 12434 15116
rect 14090 15104 14096 15156
rect 14148 15104 14154 15156
rect 14366 15104 14372 15156
rect 14424 15104 14430 15156
rect 16666 15104 16672 15156
rect 16724 15104 16730 15156
rect 17126 15104 17132 15156
rect 17184 15104 17190 15156
rect 17313 15147 17371 15153
rect 17313 15113 17325 15147
rect 17359 15144 17371 15147
rect 17770 15144 17776 15156
rect 17359 15116 17776 15144
rect 17359 15113 17371 15116
rect 17313 15107 17371 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 18509 15147 18567 15153
rect 18509 15113 18521 15147
rect 18555 15144 18567 15147
rect 18782 15144 18788 15156
rect 18555 15116 18788 15144
rect 18555 15113 18567 15116
rect 18509 15107 18567 15113
rect 18782 15104 18788 15116
rect 18840 15104 18846 15156
rect 12621 15011 12679 15017
rect 12621 15008 12633 15011
rect 12406 14980 12633 15008
rect 12621 14977 12633 14980
rect 12667 14977 12679 15011
rect 14108 15008 14136 15104
rect 15470 15036 15476 15088
rect 15528 15085 15534 15088
rect 15528 15076 15540 15085
rect 16684 15076 16712 15104
rect 18230 15076 18236 15088
rect 15528 15048 15573 15076
rect 16684 15048 18236 15076
rect 15528 15039 15540 15048
rect 15528 15036 15534 15039
rect 18230 15036 18236 15048
rect 18288 15076 18294 15088
rect 20346 15076 20352 15088
rect 18288 15048 20352 15076
rect 18288 15036 18294 15048
rect 14734 15008 14740 15020
rect 14108 14980 14740 15008
rect 12621 14971 12679 14977
rect 14734 14968 14740 14980
rect 14792 15008 14798 15020
rect 15746 15008 15752 15020
rect 14792 14980 15752 15008
rect 14792 14968 14798 14980
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 14977 17279 15011
rect 17221 14971 17279 14977
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 15008 17555 15011
rect 17589 15011 17647 15017
rect 17589 15008 17601 15011
rect 17543 14980 17601 15008
rect 17543 14977 17555 14980
rect 17497 14971 17555 14977
rect 17589 14977 17601 14980
rect 17635 14977 17647 15011
rect 17589 14971 17647 14977
rect 17236 14940 17264 14971
rect 18874 14968 18880 15020
rect 18932 15008 18938 15020
rect 19904 15017 19932 15048
rect 20346 15036 20352 15048
rect 20404 15036 20410 15088
rect 19622 15011 19680 15017
rect 19622 15008 19634 15011
rect 18932 14980 19634 15008
rect 18932 14968 18938 14980
rect 19622 14977 19634 14980
rect 19668 14977 19680 15011
rect 19622 14971 19680 14977
rect 19889 15011 19947 15017
rect 19889 14977 19901 15011
rect 19935 14977 19947 15011
rect 19889 14971 19947 14977
rect 18138 14940 18144 14952
rect 11992 14912 12388 14940
rect 17236 14912 18144 14940
rect 12253 14875 12311 14881
rect 12253 14872 12265 14875
rect 11624 14844 12265 14872
rect 11517 14835 11575 14841
rect 12253 14841 12265 14844
rect 12299 14841 12311 14875
rect 12253 14835 12311 14841
rect 11532 14804 11560 14835
rect 12360 14816 12388 14912
rect 18138 14900 18144 14912
rect 18196 14900 18202 14952
rect 16945 14875 17003 14881
rect 16945 14841 16957 14875
rect 16991 14872 17003 14875
rect 17310 14872 17316 14884
rect 16991 14844 17316 14872
rect 16991 14841 17003 14844
rect 16945 14835 17003 14841
rect 17310 14832 17316 14844
rect 17368 14832 17374 14884
rect 17773 14875 17831 14881
rect 17773 14841 17785 14875
rect 17819 14872 17831 14875
rect 17862 14872 17868 14884
rect 17819 14844 17868 14872
rect 17819 14841 17831 14844
rect 17773 14835 17831 14841
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 10980 14776 11560 14804
rect 8481 14767 8539 14773
rect 12158 14764 12164 14816
rect 12216 14764 12222 14816
rect 12342 14764 12348 14816
rect 12400 14764 12406 14816
rect 1104 14714 20792 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 10214 14714
rect 10266 14662 10278 14714
rect 10330 14662 10342 14714
rect 10394 14662 10406 14714
rect 10458 14662 10470 14714
rect 10522 14662 16214 14714
rect 16266 14662 16278 14714
rect 16330 14662 16342 14714
rect 16394 14662 16406 14714
rect 16458 14662 16470 14714
rect 16522 14662 20792 14714
rect 1104 14640 20792 14662
rect 1486 14560 1492 14612
rect 1544 14560 1550 14612
rect 2314 14560 2320 14612
rect 2372 14600 2378 14612
rect 3145 14603 3203 14609
rect 3145 14600 3157 14603
rect 2372 14572 3157 14600
rect 2372 14560 2378 14572
rect 3145 14569 3157 14572
rect 3191 14569 3203 14603
rect 3145 14563 3203 14569
rect 3694 14560 3700 14612
rect 3752 14600 3758 14612
rect 5258 14600 5264 14612
rect 3752 14572 5264 14600
rect 3752 14560 3758 14572
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 5537 14603 5595 14609
rect 5537 14569 5549 14603
rect 5583 14600 5595 14603
rect 5902 14600 5908 14612
rect 5583 14572 5908 14600
rect 5583 14569 5595 14572
rect 5537 14563 5595 14569
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 6454 14560 6460 14612
rect 6512 14560 6518 14612
rect 6730 14560 6736 14612
rect 6788 14560 6794 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 7024 14572 7481 14600
rect 1504 14464 1532 14560
rect 1673 14467 1731 14473
rect 1673 14464 1685 14467
rect 1504 14436 1685 14464
rect 1673 14433 1685 14436
rect 1719 14433 1731 14467
rect 3712 14464 3740 14560
rect 1673 14427 1731 14433
rect 2792 14436 3740 14464
rect 2792 14408 2820 14436
rect 3786 14424 3792 14476
rect 3844 14424 3850 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4706 14464 4712 14476
rect 4111 14436 4712 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 1412 14328 1440 14359
rect 2774 14356 2780 14408
rect 2832 14356 2838 14408
rect 5276 14396 5304 14560
rect 6472 14532 6500 14560
rect 6917 14535 6975 14541
rect 6917 14532 6929 14535
rect 6472 14504 6929 14532
rect 6917 14501 6929 14504
rect 6963 14501 6975 14535
rect 6917 14495 6975 14501
rect 6270 14424 6276 14476
rect 6328 14464 6334 14476
rect 7024 14464 7052 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 7469 14563 7527 14569
rect 7742 14560 7748 14612
rect 7800 14560 7806 14612
rect 8481 14603 8539 14609
rect 8481 14569 8493 14603
rect 8527 14600 8539 14603
rect 8570 14600 8576 14612
rect 8527 14572 8576 14600
rect 8527 14569 8539 14572
rect 8481 14563 8539 14569
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 11330 14560 11336 14612
rect 11388 14600 11394 14612
rect 12158 14600 12164 14612
rect 11388 14572 12164 14600
rect 11388 14560 11394 14572
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 18598 14600 18604 14612
rect 12308 14572 18604 14600
rect 12308 14560 12314 14572
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 7101 14535 7159 14541
rect 7101 14501 7113 14535
rect 7147 14532 7159 14535
rect 7147 14504 7512 14532
rect 7147 14501 7159 14504
rect 7101 14495 7159 14501
rect 6328 14436 7052 14464
rect 6328 14424 6334 14436
rect 5198 14368 5304 14396
rect 6362 14356 6368 14408
rect 6420 14396 6426 14408
rect 7484 14405 7512 14504
rect 6641 14399 6699 14405
rect 6641 14396 6653 14399
rect 6420 14368 6653 14396
rect 6420 14356 6426 14368
rect 6641 14365 6653 14368
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14365 7527 14399
rect 7469 14359 7527 14365
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14396 7711 14399
rect 7760 14396 7788 14560
rect 9646 14504 11284 14532
rect 9646 14464 9674 14504
rect 7699 14368 7788 14396
rect 8956 14436 9674 14464
rect 11256 14464 11284 14504
rect 14734 14492 14740 14544
rect 14792 14492 14798 14544
rect 12250 14464 12256 14476
rect 11256 14436 12256 14464
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 1946 14328 1952 14340
rect 1412 14300 1952 14328
rect 1946 14288 1952 14300
rect 2004 14288 2010 14340
rect 7377 14331 7435 14337
rect 7377 14328 7389 14331
rect 7024 14300 7389 14328
rect 7024 14272 7052 14300
rect 7377 14297 7389 14300
rect 7423 14297 7435 14331
rect 7484 14328 7512 14359
rect 8956 14328 8984 14436
rect 12250 14424 12256 14436
rect 12308 14424 12314 14476
rect 12342 14424 12348 14476
rect 12400 14464 12406 14476
rect 13173 14467 13231 14473
rect 13173 14464 13185 14467
rect 12400 14436 13185 14464
rect 12400 14424 12406 14436
rect 13173 14433 13185 14436
rect 13219 14433 13231 14467
rect 14752 14464 14780 14492
rect 14921 14467 14979 14473
rect 14921 14464 14933 14467
rect 14752 14436 14933 14464
rect 13173 14427 13231 14433
rect 14921 14433 14933 14436
rect 14967 14433 14979 14467
rect 14921 14427 14979 14433
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11330 14396 11336 14408
rect 11195 14368 11336 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 11425 14399 11483 14405
rect 11425 14365 11437 14399
rect 11471 14365 11483 14399
rect 11425 14359 11483 14365
rect 11440 14328 11468 14359
rect 7484 14300 8984 14328
rect 11072 14300 11468 14328
rect 11701 14331 11759 14337
rect 7377 14291 7435 14297
rect 11072 14272 11100 14300
rect 11701 14297 11713 14331
rect 11747 14297 11759 14331
rect 11701 14291 11759 14297
rect 7006 14220 7012 14272
rect 7064 14220 7070 14272
rect 11054 14220 11060 14272
rect 11112 14220 11118 14272
rect 11333 14263 11391 14269
rect 11333 14229 11345 14263
rect 11379 14260 11391 14263
rect 11716 14260 11744 14291
rect 12710 14288 12716 14340
rect 12768 14288 12774 14340
rect 15188 14331 15246 14337
rect 15188 14297 15200 14331
rect 15234 14328 15246 14331
rect 15838 14328 15844 14340
rect 15234 14300 15844 14328
rect 15234 14297 15246 14300
rect 15188 14291 15246 14297
rect 15838 14288 15844 14300
rect 15896 14288 15902 14340
rect 11379 14232 11744 14260
rect 11379 14229 11391 14232
rect 11333 14223 11391 14229
rect 15930 14220 15936 14272
rect 15988 14260 15994 14272
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 15988 14232 16313 14260
rect 15988 14220 15994 14232
rect 16301 14229 16313 14232
rect 16347 14229 16359 14263
rect 16301 14223 16359 14229
rect 16666 14220 16672 14272
rect 16724 14220 16730 14272
rect 1104 14170 20792 14192
rect 1104 14118 7214 14170
rect 7266 14118 7278 14170
rect 7330 14118 7342 14170
rect 7394 14118 7406 14170
rect 7458 14118 7470 14170
rect 7522 14118 13214 14170
rect 13266 14118 13278 14170
rect 13330 14118 13342 14170
rect 13394 14118 13406 14170
rect 13458 14118 13470 14170
rect 13522 14118 19214 14170
rect 19266 14118 19278 14170
rect 19330 14118 19342 14170
rect 19394 14118 19406 14170
rect 19458 14118 19470 14170
rect 19522 14118 20792 14170
rect 1104 14096 20792 14118
rect 2038 14016 2044 14068
rect 2096 14016 2102 14068
rect 7742 14016 7748 14068
rect 7800 14016 7806 14068
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 9125 14059 9183 14065
rect 9125 14056 9137 14059
rect 8536 14028 9137 14056
rect 8536 14016 8542 14028
rect 9125 14025 9137 14028
rect 9171 14025 9183 14059
rect 10686 14056 10692 14068
rect 9125 14019 9183 14025
rect 9232 14028 10692 14056
rect 2056 13920 2084 14016
rect 6362 13948 6368 14000
rect 6420 13988 6426 14000
rect 7101 13991 7159 13997
rect 7101 13988 7113 13991
rect 6420 13960 7113 13988
rect 6420 13948 6426 13960
rect 7101 13957 7113 13960
rect 7147 13957 7159 13991
rect 7101 13951 7159 13957
rect 6914 13929 6920 13932
rect 2225 13923 2283 13929
rect 2225 13920 2237 13923
rect 2056 13892 2237 13920
rect 2225 13889 2237 13892
rect 2271 13889 2283 13923
rect 2225 13883 2283 13889
rect 6912 13883 6920 13929
rect 6914 13880 6920 13883
rect 6972 13880 6978 13932
rect 7006 13880 7012 13932
rect 7064 13880 7070 13932
rect 7285 13923 7343 13929
rect 7285 13889 7297 13923
rect 7331 13920 7343 13923
rect 7760 13920 7788 14016
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 9232 13988 9260 14028
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 14090 14016 14096 14068
rect 14148 14016 14154 14068
rect 14369 14059 14427 14065
rect 14369 14025 14381 14059
rect 14415 14056 14427 14059
rect 14415 14028 15332 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 7892 13960 9260 13988
rect 7892 13948 7898 13960
rect 7331 13892 7788 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 8386 13880 8392 13932
rect 8444 13880 8450 13932
rect 8570 13880 8576 13932
rect 8628 13880 8634 13932
rect 8680 13929 8708 13960
rect 10134 13948 10140 14000
rect 10192 13988 10198 14000
rect 12710 13988 12716 14000
rect 10192 13960 12716 13988
rect 10192 13948 10198 13960
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 1854 13812 1860 13864
rect 1912 13852 1918 13864
rect 2133 13855 2191 13861
rect 2133 13852 2145 13855
rect 1912 13824 2145 13852
rect 1912 13812 1918 13824
rect 2133 13821 2145 13824
rect 2179 13821 2191 13855
rect 7024 13852 7052 13880
rect 8404 13852 8432 13880
rect 7024 13824 8432 13852
rect 8588 13852 8616 13880
rect 8956 13852 8984 13883
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 10045 13923 10103 13929
rect 10045 13920 10057 13923
rect 9180 13892 10057 13920
rect 9180 13880 9186 13892
rect 10045 13889 10057 13892
rect 10091 13889 10103 13923
rect 15304 13920 15332 14028
rect 16298 14016 16304 14068
rect 16356 14016 16362 14068
rect 18230 14016 18236 14068
rect 18288 14056 18294 14068
rect 18509 14059 18567 14065
rect 18509 14056 18521 14059
rect 18288 14028 18521 14056
rect 18288 14016 18294 14028
rect 18509 14025 18521 14028
rect 18555 14025 18567 14059
rect 18509 14019 18567 14025
rect 18785 14059 18843 14065
rect 18785 14025 18797 14059
rect 18831 14056 18843 14059
rect 18874 14056 18880 14068
rect 18831 14028 18880 14056
rect 18831 14025 18843 14028
rect 18785 14019 18843 14025
rect 15470 13948 15476 14000
rect 15528 13997 15534 14000
rect 15528 13991 15562 13997
rect 15550 13988 15562 13991
rect 15841 13991 15899 13997
rect 15841 13988 15853 13991
rect 15550 13960 15853 13988
rect 15550 13957 15562 13960
rect 15528 13951 15562 13957
rect 15841 13957 15853 13960
rect 15887 13957 15899 13991
rect 15841 13951 15899 13957
rect 15528 13948 15534 13951
rect 15304 13892 15884 13920
rect 10045 13883 10103 13889
rect 15856 13864 15884 13892
rect 16022 13880 16028 13932
rect 16080 13920 16086 13932
rect 16942 13929 16948 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 16080 13892 16129 13920
rect 16080 13880 16086 13892
rect 16117 13889 16129 13892
rect 16163 13920 16175 13923
rect 16925 13923 16948 13929
rect 16925 13920 16937 13923
rect 16163 13892 16937 13920
rect 16163 13889 16175 13892
rect 16117 13883 16175 13889
rect 16925 13889 16937 13892
rect 16925 13883 16948 13889
rect 16942 13880 16948 13883
rect 17000 13880 17006 13932
rect 18524 13920 18552 14019
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 19610 13948 19616 14000
rect 19668 13988 19674 14000
rect 19898 13991 19956 13997
rect 19898 13988 19910 13991
rect 19668 13960 19910 13988
rect 19668 13948 19674 13960
rect 19898 13957 19910 13960
rect 19944 13957 19956 13991
rect 19898 13951 19956 13957
rect 20165 13923 20223 13929
rect 20165 13920 20177 13923
rect 18524 13892 20177 13920
rect 20165 13889 20177 13892
rect 20211 13889 20223 13923
rect 20165 13883 20223 13889
rect 8588 13824 8984 13852
rect 2133 13815 2191 13821
rect 10502 13812 10508 13864
rect 10560 13812 10566 13864
rect 11057 13855 11115 13861
rect 11057 13821 11069 13855
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 11072 13784 11100 13815
rect 15746 13812 15752 13864
rect 15804 13812 15810 13864
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 15896 13824 15945 13852
rect 15896 13812 15902 13824
rect 15933 13821 15945 13824
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 16666 13812 16672 13864
rect 16724 13812 16730 13864
rect 10152 13756 11100 13784
rect 15764 13784 15792 13812
rect 16684 13784 16712 13812
rect 15764 13756 16712 13784
rect 6730 13676 6736 13728
rect 6788 13676 6794 13728
rect 8754 13676 8760 13728
rect 8812 13676 8818 13728
rect 9950 13676 9956 13728
rect 10008 13716 10014 13728
rect 10152 13725 10180 13756
rect 10137 13719 10195 13725
rect 10137 13716 10149 13719
rect 10008 13688 10149 13716
rect 10008 13676 10014 13688
rect 10137 13685 10149 13688
rect 10183 13685 10195 13719
rect 10137 13679 10195 13685
rect 15930 13676 15936 13728
rect 15988 13676 15994 13728
rect 18046 13676 18052 13728
rect 18104 13676 18110 13728
rect 1104 13626 20792 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 10214 13626
rect 10266 13574 10278 13626
rect 10330 13574 10342 13626
rect 10394 13574 10406 13626
rect 10458 13574 10470 13626
rect 10522 13574 16214 13626
rect 16266 13574 16278 13626
rect 16330 13574 16342 13626
rect 16394 13574 16406 13626
rect 16458 13574 16470 13626
rect 16522 13574 20792 13626
rect 1104 13552 20792 13574
rect 5064 13515 5122 13521
rect 5064 13481 5076 13515
rect 5110 13512 5122 13515
rect 6270 13512 6276 13524
rect 5110 13484 6276 13512
rect 5110 13481 5122 13484
rect 5064 13475 5122 13481
rect 6270 13472 6276 13484
rect 6328 13472 6334 13524
rect 8386 13472 8392 13524
rect 8444 13472 8450 13524
rect 11333 13515 11391 13521
rect 11333 13481 11345 13515
rect 11379 13512 11391 13515
rect 20254 13512 20260 13524
rect 11379 13484 20260 13512
rect 11379 13481 11391 13484
rect 11333 13475 11391 13481
rect 20254 13472 20260 13484
rect 20312 13472 20318 13524
rect 3142 13404 3148 13456
rect 3200 13404 3206 13456
rect 4617 13447 4675 13453
rect 4617 13413 4629 13447
rect 4663 13413 4675 13447
rect 4617 13407 4675 13413
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2038 13376 2044 13388
rect 1443 13348 2044 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2038 13336 2044 13348
rect 2096 13376 2102 13388
rect 4632 13376 4660 13407
rect 10686 13404 10692 13456
rect 10744 13444 10750 13456
rect 10744 13416 11560 13444
rect 10744 13404 10750 13416
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 2096 13348 4108 13376
rect 4632 13348 4813 13376
rect 2096 13336 2102 13348
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 3326 13308 3332 13320
rect 2832 13280 3332 13308
rect 2832 13268 2838 13280
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 4080 13317 4108 13348
rect 4801 13345 4813 13348
rect 4847 13376 4859 13379
rect 6914 13376 6920 13388
rect 4847 13348 6920 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 8754 13336 8760 13388
rect 8812 13376 8818 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8812 13348 8953 13376
rect 8812 13336 8818 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 11422 13376 11428 13388
rect 8941 13339 8999 13345
rect 10796 13348 11428 13376
rect 10796 13320 10824 13348
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4341 13311 4399 13317
rect 4341 13308 4353 13311
rect 4065 13271 4123 13277
rect 4172 13280 4353 13308
rect 1670 13200 1676 13252
rect 1728 13200 1734 13252
rect 2958 13200 2964 13252
rect 3016 13240 3022 13252
rect 3510 13240 3516 13252
rect 3016 13212 3516 13240
rect 3016 13200 3022 13212
rect 3510 13200 3516 13212
rect 3568 13240 3574 13252
rect 4172 13240 4200 13280
rect 4341 13277 4353 13280
rect 4387 13277 4399 13311
rect 4341 13271 4399 13277
rect 4485 13311 4543 13317
rect 4485 13277 4497 13311
rect 4531 13308 4543 13311
rect 4531 13277 4568 13308
rect 4485 13271 4568 13277
rect 3568 13212 4200 13240
rect 3568 13200 3574 13212
rect 4246 13200 4252 13252
rect 4304 13200 4310 13252
rect 4540 13184 4568 13271
rect 6638 13268 6644 13320
rect 6696 13268 6702 13320
rect 10778 13268 10784 13320
rect 10836 13268 10842 13320
rect 11201 13311 11259 13317
rect 11201 13277 11213 13311
rect 11247 13308 11259 13311
rect 11532 13308 11560 13416
rect 15470 13404 15476 13456
rect 15528 13404 15534 13456
rect 16942 13404 16948 13456
rect 17000 13444 17006 13456
rect 17037 13447 17095 13453
rect 17037 13444 17049 13447
rect 17000 13416 17049 13444
rect 17000 13404 17006 13416
rect 17037 13413 17049 13416
rect 17083 13413 17095 13447
rect 17037 13407 17095 13413
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13376 13231 13379
rect 13817 13379 13875 13385
rect 13817 13376 13829 13379
rect 13219 13348 13829 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 13817 13345 13829 13348
rect 13863 13376 13875 13379
rect 14090 13376 14096 13388
rect 13863 13348 14096 13376
rect 13863 13345 13875 13348
rect 13817 13339 13875 13345
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 11247 13280 11560 13308
rect 15657 13311 15715 13317
rect 11247 13277 11259 13280
rect 11201 13271 11259 13277
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 15746 13308 15752 13320
rect 15703 13280 15752 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 15930 13317 15936 13320
rect 15924 13308 15936 13317
rect 15891 13280 15936 13308
rect 15924 13271 15936 13280
rect 15930 13268 15936 13271
rect 15988 13268 15994 13320
rect 16666 13268 16672 13320
rect 16724 13308 16730 13320
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 16724 13280 17417 13308
rect 16724 13268 16730 13280
rect 17405 13277 17417 13280
rect 17451 13308 17463 13311
rect 19058 13308 19064 13320
rect 17451 13280 19064 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 5718 13200 5724 13252
rect 5776 13200 5782 13252
rect 6917 13243 6975 13249
rect 6917 13240 6929 13243
rect 6564 13212 6929 13240
rect 2314 13132 2320 13184
rect 2372 13172 2378 13184
rect 4522 13172 4528 13184
rect 2372 13144 4528 13172
rect 2372 13132 2378 13144
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 6564 13181 6592 13212
rect 6917 13209 6929 13212
rect 6963 13209 6975 13243
rect 6917 13203 6975 13209
rect 7006 13200 7012 13252
rect 7064 13240 7070 13252
rect 8665 13243 8723 13249
rect 7064 13212 7406 13240
rect 7064 13200 7070 13212
rect 8665 13209 8677 13243
rect 8711 13240 8723 13243
rect 9122 13240 9128 13252
rect 8711 13212 9128 13240
rect 8711 13209 8723 13212
rect 8665 13203 8723 13209
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 9217 13243 9275 13249
rect 9217 13209 9229 13243
rect 9263 13240 9275 13243
rect 9490 13240 9496 13252
rect 9263 13212 9496 13240
rect 9263 13209 9275 13212
rect 9217 13203 9275 13209
rect 9490 13200 9496 13212
rect 9548 13200 9554 13252
rect 10502 13240 10508 13252
rect 10442 13212 10508 13240
rect 10502 13200 10508 13212
rect 10560 13200 10566 13252
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 10965 13243 11023 13249
rect 10965 13240 10977 13243
rect 10928 13212 10977 13240
rect 10928 13200 10934 13212
rect 10965 13209 10977 13212
rect 11011 13209 11023 13243
rect 10965 13203 11023 13209
rect 11057 13243 11115 13249
rect 11057 13209 11069 13243
rect 11103 13209 11115 13243
rect 11057 13203 11115 13209
rect 14360 13243 14418 13249
rect 14360 13209 14372 13243
rect 14406 13240 14418 13243
rect 14734 13240 14740 13252
rect 14406 13212 14740 13240
rect 14406 13209 14418 13212
rect 14360 13203 14418 13209
rect 6549 13175 6607 13181
rect 6549 13141 6561 13175
rect 6595 13141 6607 13175
rect 6549 13135 6607 13141
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 9140 13172 9168 13200
rect 9582 13172 9588 13184
rect 9140 13144 9588 13172
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 11072 13172 11100 13203
rect 14734 13200 14740 13212
rect 14792 13200 14798 13252
rect 18322 13200 18328 13252
rect 18380 13240 18386 13252
rect 18794 13243 18852 13249
rect 18794 13240 18806 13243
rect 18380 13212 18806 13240
rect 18380 13200 18386 13212
rect 18794 13209 18806 13212
rect 18840 13209 18852 13243
rect 18794 13203 18852 13209
rect 10744 13144 11100 13172
rect 10744 13132 10750 13144
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 17681 13175 17739 13181
rect 17681 13172 17693 13175
rect 17460 13144 17693 13172
rect 17460 13132 17466 13144
rect 17681 13141 17693 13144
rect 17727 13141 17739 13175
rect 17681 13135 17739 13141
rect 1104 13082 20792 13104
rect 1104 13030 7214 13082
rect 7266 13030 7278 13082
rect 7330 13030 7342 13082
rect 7394 13030 7406 13082
rect 7458 13030 7470 13082
rect 7522 13030 13214 13082
rect 13266 13030 13278 13082
rect 13330 13030 13342 13082
rect 13394 13030 13406 13082
rect 13458 13030 13470 13082
rect 13522 13030 19214 13082
rect 19266 13030 19278 13082
rect 19330 13030 19342 13082
rect 19394 13030 19406 13082
rect 19458 13030 19470 13082
rect 19522 13030 20792 13082
rect 1104 13008 20792 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 2225 12971 2283 12977
rect 2225 12968 2237 12971
rect 1728 12940 2237 12968
rect 1728 12928 1734 12940
rect 2225 12937 2237 12940
rect 2271 12937 2283 12971
rect 2225 12931 2283 12937
rect 2314 12928 2320 12980
rect 2372 12928 2378 12980
rect 4341 12971 4399 12977
rect 4341 12937 4353 12971
rect 4387 12937 4399 12971
rect 4341 12931 4399 12937
rect 2332 12900 2360 12928
rect 2958 12900 2964 12912
rect 1688 12872 2360 12900
rect 2608 12872 2964 12900
rect 1688 12841 1716 12872
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 2409 12835 2467 12841
rect 2409 12832 2421 12835
rect 1673 12795 1731 12801
rect 2148 12804 2421 12832
rect 2148 12773 2176 12804
rect 2409 12801 2421 12804
rect 2455 12801 2467 12835
rect 2409 12795 2467 12801
rect 2133 12767 2191 12773
rect 2133 12733 2145 12767
rect 2179 12733 2191 12767
rect 2133 12727 2191 12733
rect 2498 12724 2504 12776
rect 2556 12764 2562 12776
rect 2608 12773 2636 12872
rect 2958 12860 2964 12872
rect 3016 12860 3022 12912
rect 3326 12860 3332 12912
rect 3384 12860 3390 12912
rect 4356 12900 4384 12931
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 4580 12940 6193 12968
rect 4580 12928 4586 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 6638 12968 6644 12980
rect 6595 12940 6644 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 9490 12928 9496 12980
rect 9548 12928 9554 12980
rect 10870 12968 10876 12980
rect 9600 12940 10876 12968
rect 4709 12903 4767 12909
rect 4709 12900 4721 12903
rect 4356 12872 4721 12900
rect 4709 12869 4721 12872
rect 4755 12869 4767 12903
rect 4709 12863 4767 12869
rect 5718 12860 5724 12912
rect 5776 12860 5782 12912
rect 8478 12900 8484 12912
rect 7024 12872 8484 12900
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12832 6515 12835
rect 6914 12832 6920 12844
rect 6503 12804 6920 12832
rect 6503 12801 6515 12804
rect 6457 12795 6515 12801
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2556 12736 2605 12764
rect 2556 12724 2562 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 2866 12724 2872 12776
rect 2924 12724 2930 12776
rect 4430 12724 4436 12776
rect 4488 12724 4494 12776
rect 7024 12708 7052 12872
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 7742 12792 7748 12844
rect 7800 12792 7806 12844
rect 9600 12841 9628 12940
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12937 11391 12971
rect 11333 12931 11391 12937
rect 11146 12900 11152 12912
rect 11086 12872 11152 12900
rect 11146 12860 11152 12872
rect 11204 12860 11210 12912
rect 11348 12900 11376 12931
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 13265 12971 13323 12977
rect 13265 12968 13277 12971
rect 11480 12940 13277 12968
rect 11480 12928 11486 12940
rect 13265 12937 13277 12940
rect 13311 12937 13323 12971
rect 13265 12931 13323 12937
rect 14734 12928 14740 12980
rect 14792 12928 14798 12980
rect 15470 12928 15476 12980
rect 15528 12968 15534 12980
rect 15749 12971 15807 12977
rect 15749 12968 15761 12971
rect 15528 12940 15761 12968
rect 15528 12928 15534 12940
rect 15749 12937 15761 12940
rect 15795 12937 15807 12971
rect 15749 12931 15807 12937
rect 15838 12928 15844 12980
rect 15896 12928 15902 12980
rect 15930 12928 15936 12980
rect 15988 12928 15994 12980
rect 17589 12971 17647 12977
rect 17589 12937 17601 12971
rect 17635 12968 17647 12971
rect 19334 12968 19340 12980
rect 17635 12940 19340 12968
rect 17635 12937 17647 12940
rect 17589 12931 17647 12937
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 11793 12903 11851 12909
rect 11793 12900 11805 12903
rect 11348 12872 11805 12900
rect 11793 12869 11805 12872
rect 11839 12869 11851 12903
rect 11793 12863 11851 12869
rect 13372 12872 14136 12900
rect 13372 12844 13400 12872
rect 14108 12844 14136 12872
rect 16022 12860 16028 12912
rect 16080 12900 16086 12912
rect 16117 12903 16175 12909
rect 16117 12900 16129 12903
rect 16080 12872 16129 12900
rect 16080 12860 16086 12872
rect 16117 12869 16129 12872
rect 16163 12869 16175 12903
rect 16117 12863 16175 12869
rect 17218 12860 17224 12912
rect 17276 12900 17282 12912
rect 17313 12903 17371 12909
rect 17313 12900 17325 12903
rect 17276 12872 17325 12900
rect 17276 12860 17282 12872
rect 17313 12869 17325 12872
rect 17359 12900 17371 12903
rect 17402 12900 17408 12912
rect 17359 12872 17408 12900
rect 17359 12869 17371 12872
rect 17313 12863 17371 12869
rect 17402 12860 17408 12872
rect 17460 12860 17466 12912
rect 18322 12900 18328 12912
rect 17512 12872 18328 12900
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12801 9643 12835
rect 9585 12795 9643 12801
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8386 12764 8392 12776
rect 8067 12736 8392 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 9858 12724 9864 12776
rect 9916 12724 9922 12776
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 2041 12699 2099 12705
rect 2041 12665 2053 12699
rect 2087 12665 2099 12699
rect 2041 12659 2099 12665
rect 2056 12628 2084 12659
rect 5718 12656 5724 12708
rect 5776 12696 5782 12708
rect 6454 12696 6460 12708
rect 5776 12668 6460 12696
rect 5776 12656 5782 12668
rect 6454 12656 6460 12668
rect 6512 12696 6518 12708
rect 7006 12696 7012 12708
rect 6512 12668 7012 12696
rect 6512 12656 6518 12668
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 2130 12628 2136 12640
rect 2056 12600 2136 12628
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10502 12628 10508 12640
rect 10008 12600 10508 12628
rect 10008 12588 10014 12600
rect 10502 12588 10508 12600
rect 10560 12628 10566 12640
rect 12912 12628 12940 12818
rect 13354 12792 13360 12844
rect 13412 12792 13418 12844
rect 13624 12835 13682 12841
rect 13624 12801 13636 12835
rect 13670 12832 13682 12835
rect 13906 12832 13912 12844
rect 13670 12804 13912 12832
rect 13670 12801 13682 12804
rect 13624 12795 13682 12801
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14090 12792 14096 12844
rect 14148 12832 14154 12844
rect 14642 12832 14648 12844
rect 14148 12804 14648 12832
rect 14148 12792 14154 12804
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12832 15531 12835
rect 15746 12832 15752 12844
rect 15519 12804 15752 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 17512 12841 17540 12872
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12832 17739 12835
rect 18046 12832 18052 12844
rect 17727 12804 18052 12832
rect 17727 12801 17739 12804
rect 17681 12795 17739 12801
rect 18046 12792 18052 12804
rect 18104 12832 18110 12844
rect 18224 12835 18282 12841
rect 18224 12832 18236 12835
rect 18104 12804 18236 12832
rect 18104 12792 18110 12804
rect 18224 12801 18236 12804
rect 18270 12832 18282 12835
rect 18966 12832 18972 12844
rect 18270 12804 18972 12832
rect 18270 12801 18282 12804
rect 18224 12795 18282 12801
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 17957 12767 18015 12773
rect 17957 12764 17969 12767
rect 17144 12736 17969 12764
rect 10560 12600 12940 12628
rect 10560 12588 10566 12600
rect 15562 12588 15568 12640
rect 15620 12588 15626 12640
rect 16942 12588 16948 12640
rect 17000 12628 17006 12640
rect 17144 12637 17172 12736
rect 17957 12733 17969 12736
rect 18003 12733 18015 12767
rect 17957 12727 18015 12733
rect 17129 12631 17187 12637
rect 17129 12628 17141 12631
rect 17000 12600 17141 12628
rect 17000 12588 17006 12600
rect 17129 12597 17141 12600
rect 17175 12597 17187 12631
rect 17129 12591 17187 12597
rect 17862 12588 17868 12640
rect 17920 12588 17926 12640
rect 1104 12538 20792 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 10214 12538
rect 10266 12486 10278 12538
rect 10330 12486 10342 12538
rect 10394 12486 10406 12538
rect 10458 12486 10470 12538
rect 10522 12486 16214 12538
rect 16266 12486 16278 12538
rect 16330 12486 16342 12538
rect 16394 12486 16406 12538
rect 16458 12486 16470 12538
rect 16522 12486 20792 12538
rect 1104 12464 20792 12486
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 2924 12396 3801 12424
rect 2924 12384 2930 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 4062 12384 4068 12436
rect 4120 12384 4126 12436
rect 4706 12384 4712 12436
rect 4764 12384 4770 12436
rect 8478 12384 8484 12436
rect 8536 12384 8542 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 9953 12427 10011 12433
rect 9953 12424 9965 12427
rect 9916 12396 9965 12424
rect 9916 12384 9922 12396
rect 9953 12393 9965 12396
rect 9999 12393 10011 12427
rect 9953 12387 10011 12393
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 11149 12427 11207 12433
rect 11149 12424 11161 12427
rect 10928 12396 11161 12424
rect 10928 12384 10934 12396
rect 11149 12393 11161 12396
rect 11195 12393 11207 12427
rect 11149 12387 11207 12393
rect 11514 12384 11520 12436
rect 11572 12384 11578 12436
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 13354 12424 13360 12436
rect 12391 12396 13360 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 3878 12356 3884 12368
rect 3252 12328 3884 12356
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 3142 12288 3148 12300
rect 2179 12260 3148 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 3252 12232 3280 12328
rect 3878 12316 3884 12328
rect 3936 12316 3942 12368
rect 3605 12291 3663 12297
rect 3605 12257 3617 12291
rect 3651 12288 3663 12291
rect 4080 12288 4108 12384
rect 10778 12288 10784 12300
rect 3651 12260 4108 12288
rect 3651 12257 3663 12260
rect 3605 12251 3663 12257
rect 1854 12180 1860 12232
rect 1912 12180 1918 12232
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4080 12220 4108 12260
rect 8496 12260 10784 12288
rect 4019 12192 4108 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 2130 12112 2136 12164
rect 2188 12112 2194 12164
rect 2148 12084 2176 12112
rect 3804 12084 3832 12183
rect 4522 12180 4528 12232
rect 4580 12220 4586 12232
rect 8496 12229 8524 12260
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 4801 12223 4859 12229
rect 4801 12220 4813 12223
rect 4580 12192 4813 12220
rect 4580 12180 4586 12192
rect 4801 12189 4813 12192
rect 4847 12220 4859 12223
rect 8297 12223 8355 12229
rect 4847 12192 5488 12220
rect 4847 12189 4859 12192
rect 4801 12183 4859 12189
rect 5460 12096 5488 12192
rect 8297 12189 8309 12223
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 8481 12183 8539 12189
rect 8772 12192 8953 12220
rect 8312 12152 8340 12183
rect 8772 12152 8800 12192
rect 8941 12189 8953 12192
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 9033 12223 9091 12229
rect 9033 12189 9045 12223
rect 9079 12220 9091 12223
rect 9490 12220 9496 12232
rect 9079 12192 9496 12220
rect 9079 12189 9091 12192
rect 9033 12183 9091 12189
rect 9490 12180 9496 12192
rect 9548 12220 9554 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9548 12192 9781 12220
rect 9548 12180 9554 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12220 10011 12223
rect 10686 12220 10692 12232
rect 9999 12192 10692 12220
rect 9999 12189 10011 12192
rect 9953 12183 10011 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10888 12229 10916 12384
rect 10965 12359 11023 12365
rect 10965 12325 10977 12359
rect 11011 12356 11023 12359
rect 11532 12356 11560 12384
rect 11011 12328 11560 12356
rect 11011 12325 11023 12328
rect 10965 12319 11023 12325
rect 12452 12232 12480 12396
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 13817 12427 13875 12433
rect 13817 12393 13829 12427
rect 13863 12424 13875 12427
rect 13906 12424 13912 12436
rect 13863 12396 13912 12424
rect 13863 12393 13875 12396
rect 13817 12387 13875 12393
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 14645 12427 14703 12433
rect 14645 12393 14657 12427
rect 14691 12424 14703 12427
rect 16025 12427 16083 12433
rect 16025 12424 16037 12427
rect 14691 12396 16037 12424
rect 14691 12393 14703 12396
rect 14645 12387 14703 12393
rect 16025 12393 16037 12396
rect 16071 12393 16083 12427
rect 16025 12387 16083 12393
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11296 12192 11345 12220
rect 11296 12180 11302 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 12434 12180 12440 12232
rect 12492 12180 12498 12232
rect 13924 12220 13952 12384
rect 14090 12316 14096 12368
rect 14148 12356 14154 12368
rect 14734 12356 14740 12368
rect 14148 12328 14740 12356
rect 14148 12316 14154 12328
rect 14734 12316 14740 12328
rect 14792 12316 14798 12368
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 16316 12356 16344 12387
rect 18322 12384 18328 12436
rect 18380 12424 18386 12436
rect 18874 12424 18880 12436
rect 18380 12396 18880 12424
rect 18380 12384 18386 12396
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 15252 12328 16344 12356
rect 15252 12316 15258 12328
rect 16942 12248 16948 12300
rect 17000 12248 17006 12300
rect 18877 12291 18935 12297
rect 18877 12257 18889 12291
rect 18923 12288 18935 12291
rect 19334 12288 19340 12300
rect 18923 12260 19340 12288
rect 18923 12257 18935 12260
rect 18877 12251 18935 12257
rect 19334 12248 19340 12260
rect 19392 12288 19398 12300
rect 19392 12260 19656 12288
rect 19392 12248 19398 12260
rect 19628 12232 19656 12260
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13924 12192 14289 12220
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 15562 12180 15568 12232
rect 15620 12220 15626 12232
rect 15620 12192 15976 12220
rect 15620 12180 15626 12192
rect 12682 12155 12740 12161
rect 12682 12152 12694 12155
rect 8312 12124 8800 12152
rect 8772 12096 8800 12124
rect 12544 12124 12694 12152
rect 12544 12096 12572 12124
rect 12682 12121 12694 12124
rect 12728 12121 12740 12155
rect 12682 12115 12740 12121
rect 15838 12112 15844 12164
rect 15896 12112 15902 12164
rect 15948 12152 15976 12192
rect 16298 12180 16304 12232
rect 16356 12180 16362 12232
rect 16390 12180 16396 12232
rect 16448 12180 16454 12232
rect 17218 12229 17224 12232
rect 17212 12183 17224 12229
rect 17276 12220 17282 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 17276 12192 18705 12220
rect 17218 12180 17224 12183
rect 17276 12180 17282 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 18966 12180 18972 12232
rect 19024 12180 19030 12232
rect 19610 12180 19616 12232
rect 19668 12180 19674 12232
rect 16041 12155 16099 12161
rect 16041 12152 16053 12155
rect 15948 12124 16053 12152
rect 16041 12121 16053 12124
rect 16087 12121 16099 12155
rect 16041 12115 16099 12121
rect 2148 12056 3832 12084
rect 5442 12044 5448 12096
rect 5500 12044 5506 12096
rect 8754 12044 8760 12096
rect 8812 12044 8818 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 12584 12056 14381 12084
rect 12584 12044 12590 12056
rect 14369 12053 14381 12056
rect 14415 12053 14427 12087
rect 14369 12047 14427 12053
rect 14458 12044 14464 12096
rect 14516 12044 14522 12096
rect 16206 12044 16212 12096
rect 16264 12044 16270 12096
rect 16666 12044 16672 12096
rect 16724 12044 16730 12096
rect 18322 12044 18328 12096
rect 18380 12044 18386 12096
rect 18506 12044 18512 12096
rect 18564 12044 18570 12096
rect 1104 11994 20792 12016
rect 1104 11942 7214 11994
rect 7266 11942 7278 11994
rect 7330 11942 7342 11994
rect 7394 11942 7406 11994
rect 7458 11942 7470 11994
rect 7522 11942 13214 11994
rect 13266 11942 13278 11994
rect 13330 11942 13342 11994
rect 13394 11942 13406 11994
rect 13458 11942 13470 11994
rect 13522 11942 19214 11994
rect 19266 11942 19278 11994
rect 19330 11942 19342 11994
rect 19394 11942 19406 11994
rect 19458 11942 19470 11994
rect 19522 11942 20792 11994
rect 1104 11920 20792 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2130 11880 2136 11892
rect 1627 11852 2136 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 2498 11840 2504 11892
rect 2556 11840 2562 11892
rect 4341 11883 4399 11889
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 4522 11880 4528 11892
rect 4387 11852 4528 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 14277 11883 14335 11889
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 15194 11880 15200 11892
rect 14323 11852 15200 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 15673 11883 15731 11889
rect 15673 11880 15685 11883
rect 15620 11852 15685 11880
rect 15620 11840 15626 11852
rect 15673 11849 15685 11852
rect 15719 11880 15731 11883
rect 15719 11852 15792 11880
rect 15719 11849 15731 11852
rect 15673 11843 15731 11849
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 14458 11812 14464 11824
rect 13872 11784 14464 11812
rect 13872 11772 13878 11784
rect 14458 11772 14464 11784
rect 14516 11772 14522 11824
rect 15286 11772 15292 11824
rect 15344 11812 15350 11824
rect 15473 11815 15531 11821
rect 15473 11812 15485 11815
rect 15344 11784 15485 11812
rect 15344 11772 15350 11784
rect 15473 11781 15485 11784
rect 15519 11781 15531 11815
rect 15473 11775 15531 11781
rect 1394 11704 1400 11756
rect 1452 11704 1458 11756
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 14001 11747 14059 11753
rect 14001 11744 14013 11747
rect 12584 11716 14013 11744
rect 12584 11704 12590 11716
rect 14001 11713 14013 11716
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 14090 11704 14096 11756
rect 14148 11704 14154 11756
rect 15488 11676 15516 11775
rect 15764 11744 15792 11852
rect 15838 11840 15844 11892
rect 15896 11840 15902 11892
rect 16206 11840 16212 11892
rect 16264 11840 16270 11892
rect 16301 11883 16359 11889
rect 16301 11849 16313 11883
rect 16347 11880 16359 11883
rect 16390 11880 16396 11892
rect 16347 11852 16396 11880
rect 16347 11849 16359 11852
rect 16301 11843 16359 11849
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 16666 11840 16672 11892
rect 16724 11880 16730 11892
rect 18141 11883 18199 11889
rect 16724 11852 18092 11880
rect 16724 11840 16730 11852
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15764 11716 15945 11744
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16025 11679 16083 11685
rect 16025 11676 16037 11679
rect 15488 11648 16037 11676
rect 16025 11645 16037 11648
rect 16071 11645 16083 11679
rect 16224 11676 16252 11840
rect 16942 11772 16948 11824
rect 17000 11772 17006 11824
rect 17310 11772 17316 11824
rect 17368 11772 17374 11824
rect 18064 11821 18092 11852
rect 18141 11849 18153 11883
rect 18187 11849 18199 11883
rect 18141 11843 18199 11849
rect 18049 11815 18107 11821
rect 18049 11781 18061 11815
rect 18095 11781 18107 11815
rect 18049 11775 18107 11781
rect 17497 11747 17555 11753
rect 17497 11713 17509 11747
rect 17543 11744 17555 11747
rect 18156 11744 18184 11843
rect 18506 11840 18512 11892
rect 18564 11840 18570 11892
rect 18874 11840 18880 11892
rect 18932 11840 18938 11892
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 20070 11880 20076 11892
rect 19116 11852 20076 11880
rect 19116 11840 19122 11852
rect 20070 11840 20076 11852
rect 20128 11880 20134 11892
rect 20128 11852 20300 11880
rect 20128 11840 20134 11852
rect 18524 11812 18552 11840
rect 17543 11716 18184 11744
rect 18248 11784 18552 11812
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 17589 11679 17647 11685
rect 17589 11676 17601 11679
rect 16224 11648 17601 11676
rect 16025 11639 16083 11645
rect 17589 11645 17601 11648
rect 17635 11645 17647 11679
rect 17589 11639 17647 11645
rect 17770 11636 17776 11688
rect 17828 11636 17834 11688
rect 18248 11685 18276 11784
rect 19610 11772 19616 11824
rect 19668 11812 19674 11824
rect 19990 11815 20048 11821
rect 19990 11812 20002 11815
rect 19668 11784 20002 11812
rect 19668 11772 19674 11784
rect 19990 11781 20002 11784
rect 20036 11781 20048 11815
rect 19990 11775 20048 11781
rect 18322 11704 18328 11756
rect 18380 11704 18386 11756
rect 20272 11753 20300 11852
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11713 20315 11747
rect 20257 11707 20315 11713
rect 17865 11679 17923 11685
rect 17865 11645 17877 11679
rect 17911 11645 17923 11679
rect 17865 11639 17923 11645
rect 17957 11679 18015 11685
rect 17957 11645 17969 11679
rect 18003 11676 18015 11679
rect 18233 11679 18291 11685
rect 18003 11648 18184 11676
rect 18003 11645 18015 11648
rect 17957 11639 18015 11645
rect 13906 11500 13912 11552
rect 13964 11500 13970 11552
rect 15657 11543 15715 11549
rect 15657 11509 15669 11543
rect 15703 11540 15715 11543
rect 16114 11540 16120 11552
rect 15703 11512 16120 11540
rect 15703 11509 15715 11512
rect 15657 11503 15715 11509
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 17880 11540 17908 11639
rect 18156 11608 18184 11648
rect 18233 11645 18245 11679
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11676 18475 11679
rect 18874 11676 18880 11688
rect 18463 11648 18880 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 18432 11608 18460 11639
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 18156 11580 18460 11608
rect 18322 11540 18328 11552
rect 17880 11512 18328 11540
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 1104 11450 20792 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 10214 11450
rect 10266 11398 10278 11450
rect 10330 11398 10342 11450
rect 10394 11398 10406 11450
rect 10458 11398 10470 11450
rect 10522 11398 16214 11450
rect 16266 11398 16278 11450
rect 16330 11398 16342 11450
rect 16394 11398 16406 11450
rect 16458 11398 16470 11450
rect 16522 11398 20792 11450
rect 1104 11376 20792 11398
rect 9125 11339 9183 11345
rect 3252 11308 5764 11336
rect 3252 11280 3280 11308
rect 3234 11228 3240 11280
rect 3292 11228 3298 11280
rect 2774 11200 2780 11212
rect 1596 11172 2780 11200
rect 1596 11141 1624 11172
rect 2774 11160 2780 11172
rect 2832 11160 2838 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 5442 11200 5448 11212
rect 4479 11172 5448 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 2271 11104 2329 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 2866 11092 2872 11144
rect 2924 11092 2930 11144
rect 5736 11132 5764 11308
rect 9125 11305 9137 11339
rect 9171 11336 9183 11339
rect 9214 11336 9220 11348
rect 9171 11308 9220 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 9582 11296 9588 11348
rect 9640 11296 9646 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11514 11336 11520 11348
rect 11112 11308 11520 11336
rect 11112 11296 11118 11308
rect 11514 11296 11520 11308
rect 11572 11336 11578 11348
rect 11885 11339 11943 11345
rect 11885 11336 11897 11339
rect 11572 11308 11897 11336
rect 11572 11296 11578 11308
rect 11885 11305 11897 11308
rect 11931 11305 11943 11339
rect 11885 11299 11943 11305
rect 12345 11339 12403 11345
rect 12345 11305 12357 11339
rect 12391 11336 12403 11339
rect 12434 11336 12440 11348
rect 12391 11308 12440 11336
rect 12391 11305 12403 11308
rect 12345 11299 12403 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 12526 11296 12532 11348
rect 12584 11296 12590 11348
rect 9309 11271 9367 11277
rect 9309 11237 9321 11271
rect 9355 11237 9367 11271
rect 9309 11231 9367 11237
rect 9677 11271 9735 11277
rect 9677 11237 9689 11271
rect 9723 11268 9735 11271
rect 9723 11240 11468 11268
rect 9723 11237 9735 11240
rect 9677 11231 9735 11237
rect 6273 11135 6331 11141
rect 6273 11132 6285 11135
rect 5736 11104 6285 11132
rect 6273 11101 6285 11104
rect 6319 11101 6331 11135
rect 6273 11095 6331 11101
rect 8478 11092 8484 11144
rect 8536 11092 8542 11144
rect 9324 11132 9352 11231
rect 10042 11160 10048 11212
rect 10100 11200 10106 11212
rect 10229 11203 10287 11209
rect 10229 11200 10241 11203
rect 10100 11172 10241 11200
rect 10100 11160 10106 11172
rect 10229 11169 10241 11172
rect 10275 11169 10287 11203
rect 10229 11163 10287 11169
rect 10870 11160 10876 11212
rect 10928 11160 10934 11212
rect 11330 11160 11336 11212
rect 11388 11160 11394 11212
rect 9401 11135 9459 11141
rect 9401 11132 9413 11135
rect 9324 11104 9413 11132
rect 9401 11101 9413 11104
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 10888 11132 10916 11160
rect 10735 11104 10916 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 3970 11024 3976 11076
rect 4028 11024 4034 11076
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 4614 11064 4620 11076
rect 4203 11036 4620 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 4706 11024 4712 11076
rect 4764 11024 4770 11076
rect 6641 11067 6699 11073
rect 6641 11033 6653 11067
rect 6687 11064 6699 11067
rect 8386 11064 8392 11076
rect 6687 11036 8392 11064
rect 6687 11033 6699 11036
rect 6641 11027 6699 11033
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 8941 11067 8999 11073
rect 8941 11064 8953 11067
rect 8720 11036 8953 11064
rect 8720 11024 8726 11036
rect 8941 11033 8953 11036
rect 8987 11033 8999 11067
rect 9141 11067 9199 11073
rect 9141 11064 9153 11067
rect 8941 11027 8999 11033
rect 9048 11036 9153 11064
rect 9048 11008 9076 11036
rect 9141 11033 9153 11036
rect 9187 11033 9199 11067
rect 9141 11027 9199 11033
rect 9858 11024 9864 11076
rect 9916 11024 9922 11076
rect 10045 11067 10103 11073
rect 10045 11033 10057 11067
rect 10091 11064 10103 11067
rect 10428 11064 10456 11095
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 11440 11141 11468 11240
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 16942 11200 16948 11212
rect 16715 11172 16948 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 16942 11160 16948 11172
rect 17000 11200 17006 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 17000 11172 18613 11200
rect 17000 11160 17006 11172
rect 18601 11169 18613 11172
rect 18647 11200 18659 11203
rect 18969 11203 19027 11209
rect 18969 11200 18981 11203
rect 18647 11172 18981 11200
rect 18647 11169 18659 11172
rect 18601 11163 18659 11169
rect 18969 11169 18981 11172
rect 19015 11169 19027 11203
rect 18969 11163 19027 11169
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 13653 11135 13711 11141
rect 13653 11101 13665 11135
rect 13699 11132 13711 11135
rect 13814 11132 13820 11144
rect 13699 11104 13820 11132
rect 13699 11101 13711 11104
rect 13653 11095 13711 11101
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 13909 11135 13967 11141
rect 13909 11101 13921 11135
rect 13955 11132 13967 11135
rect 14642 11132 14648 11144
rect 13955 11104 14648 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 14642 11092 14648 11104
rect 14700 11132 14706 11144
rect 14700 11104 14780 11132
rect 14700 11092 14706 11104
rect 10091 11036 10456 11064
rect 10597 11067 10655 11073
rect 10091 11033 10103 11036
rect 10045 11027 10103 11033
rect 10597 11033 10609 11067
rect 10643 11064 10655 11067
rect 10980 11064 11008 11092
rect 10643 11036 11008 11064
rect 10643 11033 10655 11036
rect 10597 11027 10655 11033
rect 2314 10956 2320 11008
rect 2372 10996 2378 11008
rect 2501 10999 2559 11005
rect 2501 10996 2513 10999
rect 2372 10968 2513 10996
rect 2372 10956 2378 10968
rect 2501 10965 2513 10968
rect 2547 10965 2559 10999
rect 2501 10959 2559 10965
rect 2682 10956 2688 11008
rect 2740 10956 2746 11008
rect 4341 10999 4399 11005
rect 4341 10965 4353 10999
rect 4387 10996 4399 10999
rect 4522 10996 4528 11008
rect 4387 10968 4528 10996
rect 4387 10965 4399 10968
rect 4341 10959 4399 10965
rect 4522 10956 4528 10968
rect 4580 10996 4586 11008
rect 5350 10996 5356 11008
rect 4580 10968 5356 10996
rect 4580 10956 4586 10968
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 5718 10956 5724 11008
rect 5776 10996 5782 11008
rect 6181 10999 6239 11005
rect 6181 10996 6193 10999
rect 5776 10968 6193 10996
rect 5776 10956 5782 10968
rect 6181 10965 6193 10968
rect 6227 10965 6239 10999
rect 6181 10959 6239 10965
rect 8294 10956 8300 11008
rect 8352 10956 8358 11008
rect 9030 10956 9036 11008
rect 9088 10956 9094 11008
rect 11606 10956 11612 11008
rect 11664 10956 11670 11008
rect 14752 11005 14780 11104
rect 16114 11024 16120 11076
rect 16172 11064 16178 11076
rect 16298 11064 16304 11076
rect 16172 11036 16304 11064
rect 16172 11024 16178 11036
rect 16298 11024 16304 11036
rect 16356 11064 16362 11076
rect 16402 11067 16460 11073
rect 16402 11064 16414 11067
rect 16356 11036 16414 11064
rect 16356 11024 16362 11036
rect 16402 11033 16414 11036
rect 16448 11033 16460 11067
rect 16402 11027 16460 11033
rect 14737 10999 14795 11005
rect 14737 10965 14749 10999
rect 14783 10996 14795 10999
rect 15010 10996 15016 11008
rect 14783 10968 15016 10996
rect 14783 10965 14795 10968
rect 14737 10959 14795 10965
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 15286 10956 15292 11008
rect 15344 10956 15350 11008
rect 1104 10906 20792 10928
rect 1104 10854 7214 10906
rect 7266 10854 7278 10906
rect 7330 10854 7342 10906
rect 7394 10854 7406 10906
rect 7458 10854 7470 10906
rect 7522 10854 13214 10906
rect 13266 10854 13278 10906
rect 13330 10854 13342 10906
rect 13394 10854 13406 10906
rect 13458 10854 13470 10906
rect 13522 10854 19214 10906
rect 19266 10854 19278 10906
rect 19330 10854 19342 10906
rect 19394 10854 19406 10906
rect 19458 10854 19470 10906
rect 19522 10854 20792 10906
rect 1104 10832 20792 10854
rect 2314 10792 2320 10804
rect 2240 10764 2320 10792
rect 2240 10665 2268 10764
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 4028 10764 4077 10792
rect 4028 10752 4034 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 4065 10755 4123 10761
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 4764 10764 5181 10792
rect 4764 10752 4770 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5316 10764 6408 10792
rect 5316 10752 5322 10764
rect 2498 10724 2504 10736
rect 2332 10696 2504 10724
rect 2332 10665 2360 10696
rect 2498 10684 2504 10696
rect 2556 10684 2562 10736
rect 3234 10684 3240 10736
rect 3292 10684 3298 10736
rect 4985 10727 5043 10733
rect 4985 10724 4997 10727
rect 4356 10696 4997 10724
rect 4356 10665 4384 10696
rect 4985 10693 4997 10696
rect 5031 10724 5043 10727
rect 5031 10696 5396 10724
rect 5031 10693 5043 10696
rect 4985 10687 5043 10693
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 4341 10659 4399 10665
rect 4341 10625 4353 10659
rect 4387 10625 4399 10659
rect 4341 10619 4399 10625
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10625 4491 10659
rect 4433 10619 4491 10625
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 4157 10591 4215 10597
rect 4157 10588 4169 10591
rect 2639 10560 4169 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 4157 10557 4169 10560
rect 4203 10557 4215 10591
rect 4448 10588 4476 10619
rect 4522 10616 4528 10668
rect 4580 10616 4586 10668
rect 5368 10665 5396 10696
rect 5718 10684 5724 10736
rect 5776 10684 5782 10736
rect 6380 10665 6408 10764
rect 9214 10752 9220 10804
rect 9272 10792 9278 10804
rect 9447 10795 9505 10801
rect 9447 10792 9459 10795
rect 9272 10764 9459 10792
rect 9272 10752 9278 10764
rect 9447 10761 9459 10764
rect 9493 10761 9505 10795
rect 9447 10755 9505 10761
rect 9858 10752 9864 10804
rect 9916 10752 9922 10804
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10870 10792 10876 10804
rect 10091 10764 10876 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 11146 10752 11152 10804
rect 11204 10752 11210 10804
rect 12158 10792 12164 10804
rect 11256 10764 12164 10792
rect 6472 10696 6960 10724
rect 4643 10659 4701 10665
rect 4643 10656 4655 10659
rect 4632 10625 4655 10656
rect 4689 10625 4701 10659
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4632 10619 4701 10625
rect 4816 10628 4905 10656
rect 4157 10551 4215 10557
rect 4356 10560 4476 10588
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4356 10452 4384 10560
rect 4632 10532 4660 10619
rect 4816 10600 4844 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5445 10659 5503 10665
rect 5445 10625 5457 10659
rect 5491 10656 5503 10659
rect 6181 10659 6239 10665
rect 5491 10628 5948 10656
rect 5491 10625 5503 10628
rect 5445 10619 5503 10625
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 4614 10480 4620 10532
rect 4672 10480 4678 10532
rect 5092 10520 5120 10619
rect 4724 10492 5120 10520
rect 4724 10464 4752 10492
rect 5460 10464 5488 10619
rect 5920 10597 5948 10628
rect 6181 10625 6193 10659
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6365 10659 6423 10665
rect 6365 10625 6377 10659
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 6196 10588 6224 10619
rect 6472 10588 6500 10696
rect 6546 10616 6552 10668
rect 6604 10616 6610 10668
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 6196 10560 6500 10588
rect 5905 10551 5963 10557
rect 5828 10520 5856 10551
rect 5997 10523 6055 10529
rect 5997 10520 6009 10523
rect 5828 10492 6009 10520
rect 5997 10489 6009 10492
rect 6043 10520 6055 10523
rect 6748 10520 6776 10619
rect 6932 10600 6960 10696
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 11256 10724 11284 10764
rect 12158 10752 12164 10764
rect 12216 10792 12222 10804
rect 12710 10792 12716 10804
rect 12216 10764 12716 10792
rect 12216 10752 12222 10764
rect 12710 10752 12716 10764
rect 12768 10792 12774 10804
rect 13449 10795 13507 10801
rect 12768 10764 12940 10792
rect 12768 10752 12774 10764
rect 9088 10696 11284 10724
rect 9088 10684 9094 10696
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 11793 10727 11851 10733
rect 11793 10724 11805 10727
rect 11388 10696 11805 10724
rect 11388 10684 11394 10696
rect 11793 10693 11805 10696
rect 11839 10693 11851 10727
rect 11793 10687 11851 10693
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7742 10656 7748 10668
rect 7607 10628 7748 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 7668 10597 7696 10628
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 11514 10616 11520 10668
rect 11572 10616 11578 10668
rect 12912 10642 12940 10764
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 13814 10792 13820 10804
rect 13495 10764 13820 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 16298 10752 16304 10804
rect 16356 10752 16362 10804
rect 16942 10752 16948 10804
rect 17000 10752 17006 10804
rect 18417 10795 18475 10801
rect 18417 10761 18429 10795
rect 18463 10761 18475 10795
rect 18417 10755 18475 10761
rect 14584 10727 14642 10733
rect 14584 10693 14596 10727
rect 14630 10724 14642 10727
rect 15286 10724 15292 10736
rect 14630 10696 15292 10724
rect 14630 10693 14642 10696
rect 14584 10687 14642 10693
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 14829 10659 14887 10665
rect 14829 10625 14841 10659
rect 14875 10656 14887 10659
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14875 10628 14933 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 14921 10625 14933 10628
rect 14967 10656 14979 10659
rect 15010 10656 15016 10668
rect 14967 10628 15016 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 15188 10659 15246 10665
rect 15188 10625 15200 10659
rect 15234 10656 15246 10659
rect 15470 10656 15476 10668
rect 15234 10628 15476 10656
rect 15234 10625 15246 10628
rect 15188 10619 15246 10625
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 16960 10656 16988 10752
rect 18432 10724 18460 10755
rect 18506 10724 18512 10736
rect 18432 10696 18512 10724
rect 18506 10684 18512 10696
rect 18564 10724 18570 10736
rect 19806 10727 19864 10733
rect 19806 10724 19818 10727
rect 18564 10696 19818 10724
rect 18564 10684 18570 10696
rect 19806 10693 19818 10696
rect 19852 10693 19864 10727
rect 19806 10687 19864 10693
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16960 10628 17049 10656
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 17304 10659 17362 10665
rect 17304 10625 17316 10659
rect 17350 10656 17362 10659
rect 18230 10656 18236 10668
rect 17350 10628 18236 10656
rect 17350 10625 17362 10628
rect 17304 10619 17362 10625
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 20070 10616 20076 10668
rect 20128 10616 20134 10668
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 8021 10591 8079 10597
rect 7699 10560 7733 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 8021 10557 8033 10591
rect 8067 10588 8079 10591
rect 8294 10588 8300 10600
rect 8067 10560 8300 10588
rect 8067 10557 8079 10560
rect 8021 10551 8079 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 10042 10548 10048 10600
rect 10100 10548 10106 10600
rect 10134 10548 10140 10600
rect 10192 10588 10198 10600
rect 10502 10588 10508 10600
rect 10192 10560 10508 10588
rect 10192 10548 10198 10560
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 13265 10591 13323 10597
rect 13265 10588 13277 10591
rect 11020 10560 13277 10588
rect 11020 10548 11026 10560
rect 13265 10557 13277 10560
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 6043 10492 6776 10520
rect 10060 10520 10088 10548
rect 10413 10523 10471 10529
rect 10413 10520 10425 10523
rect 10060 10492 10425 10520
rect 6043 10489 6055 10492
rect 5997 10483 6055 10489
rect 10413 10489 10425 10492
rect 10459 10489 10471 10523
rect 10413 10483 10471 10489
rect 4120 10424 4384 10452
rect 4120 10412 4126 10424
rect 4706 10412 4712 10464
rect 4764 10412 4770 10464
rect 5442 10412 5448 10464
rect 5500 10412 5506 10464
rect 6089 10455 6147 10461
rect 6089 10421 6101 10455
rect 6135 10452 6147 10455
rect 6730 10452 6736 10464
rect 6135 10424 6736 10452
rect 6135 10421 6147 10424
rect 6089 10415 6147 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 6917 10455 6975 10461
rect 6917 10421 6929 10455
rect 6963 10452 6975 10455
rect 7374 10452 7380 10464
rect 6963 10424 7380 10452
rect 6963 10421 6975 10424
rect 6917 10415 6975 10421
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 10980 10452 11008 10548
rect 10091 10424 11008 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 18322 10412 18328 10464
rect 18380 10452 18386 10464
rect 18693 10455 18751 10461
rect 18693 10452 18705 10455
rect 18380 10424 18705 10452
rect 18380 10412 18386 10424
rect 18693 10421 18705 10424
rect 18739 10421 18751 10455
rect 18693 10415 18751 10421
rect 1104 10362 20792 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 10214 10362
rect 10266 10310 10278 10362
rect 10330 10310 10342 10362
rect 10394 10310 10406 10362
rect 10458 10310 10470 10362
rect 10522 10310 16214 10362
rect 16266 10310 16278 10362
rect 16330 10310 16342 10362
rect 16394 10310 16406 10362
rect 16458 10310 16470 10362
rect 16522 10310 20792 10362
rect 1104 10288 20792 10310
rect 1578 10208 1584 10260
rect 1636 10208 1642 10260
rect 2120 10251 2178 10257
rect 2120 10217 2132 10251
rect 2166 10248 2178 10251
rect 2682 10248 2688 10260
rect 2166 10220 2688 10248
rect 2166 10217 2178 10220
rect 2120 10211 2178 10217
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 2866 10208 2872 10260
rect 2924 10248 2930 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 2924 10220 3801 10248
rect 2924 10208 2930 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4798 10248 4804 10260
rect 4028 10220 4804 10248
rect 4028 10208 4034 10220
rect 4798 10208 4804 10220
rect 4856 10248 4862 10260
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 4856 10220 4905 10248
rect 4856 10208 4862 10220
rect 4893 10217 4905 10220
rect 4939 10217 4951 10251
rect 4893 10211 4951 10217
rect 5077 10251 5135 10257
rect 5077 10217 5089 10251
rect 5123 10248 5135 10251
rect 5258 10248 5264 10260
rect 5123 10220 5264 10248
rect 5123 10217 5135 10220
rect 5077 10211 5135 10217
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5537 10251 5595 10257
rect 5537 10248 5549 10251
rect 5500 10220 5549 10248
rect 5500 10208 5506 10220
rect 5537 10217 5549 10220
rect 5583 10217 5595 10251
rect 5537 10211 5595 10217
rect 5718 10208 5724 10260
rect 5776 10208 5782 10260
rect 5905 10251 5963 10257
rect 5905 10217 5917 10251
rect 5951 10248 5963 10251
rect 6089 10251 6147 10257
rect 5951 10220 6040 10248
rect 5951 10217 5963 10220
rect 5905 10211 5963 10217
rect 1596 10053 1624 10208
rect 5736 10180 5764 10208
rect 6012 10180 6040 10220
rect 6089 10217 6101 10251
rect 6135 10248 6147 10251
rect 8389 10251 8447 10257
rect 6135 10220 7972 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 6273 10183 6331 10189
rect 6273 10180 6285 10183
rect 4264 10152 4660 10180
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 2498 10112 2504 10124
rect 1903 10084 2504 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10013 1639 10047
rect 1581 10007 1639 10013
rect 3234 10004 3240 10056
rect 3292 10004 3298 10056
rect 4264 10053 4292 10152
rect 4632 10124 4660 10152
rect 5092 10152 5948 10180
rect 6012 10152 6285 10180
rect 4341 10115 4399 10121
rect 4341 10081 4353 10115
rect 4387 10081 4399 10115
rect 4341 10075 4399 10081
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4356 9976 4384 10075
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 4798 10112 4804 10124
rect 4672 10084 4804 10112
rect 4672 10072 4678 10084
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 4706 9976 4712 9988
rect 3620 9948 4712 9976
rect 1670 9868 1676 9920
rect 1728 9868 1734 9920
rect 3620 9917 3648 9948
rect 4706 9936 4712 9948
rect 4764 9936 4770 9988
rect 4925 9979 4983 9985
rect 4925 9945 4937 9979
rect 4971 9976 4983 9979
rect 5092 9976 5120 10152
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5408 10084 5672 10112
rect 5408 10072 5414 10084
rect 5644 10053 5672 10084
rect 5718 10072 5724 10124
rect 5776 10072 5782 10124
rect 5920 10053 5948 10152
rect 6273 10149 6285 10152
rect 6319 10180 6331 10183
rect 6362 10180 6368 10192
rect 6319 10152 6368 10180
rect 6319 10149 6331 10152
rect 6273 10143 6331 10149
rect 6362 10140 6368 10152
rect 6420 10180 6426 10192
rect 6638 10180 6644 10192
rect 6420 10152 6644 10180
rect 6420 10140 6426 10152
rect 6638 10140 6644 10152
rect 6696 10140 6702 10192
rect 7944 10180 7972 10220
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 8478 10248 8484 10260
rect 8435 10220 8484 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 9490 10208 9496 10260
rect 9548 10208 9554 10260
rect 15470 10208 15476 10260
rect 15528 10208 15534 10260
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16942 10248 16948 10260
rect 16531 10220 16948 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 9309 10183 9367 10189
rect 9309 10180 9321 10183
rect 7944 10152 9321 10180
rect 9309 10149 9321 10152
rect 9355 10149 9367 10183
rect 9309 10143 9367 10149
rect 7374 10072 7380 10124
rect 7432 10112 7438 10124
rect 7745 10115 7803 10121
rect 7745 10112 7757 10115
rect 7432 10084 7757 10112
rect 7432 10072 7438 10084
rect 7745 10081 7757 10084
rect 7791 10081 7803 10115
rect 7745 10075 7803 10081
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9824 10084 10057 10112
rect 9824 10072 9830 10084
rect 10045 10081 10057 10084
rect 10091 10112 10103 10115
rect 11514 10112 11520 10124
rect 10091 10084 11520 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 11514 10072 11520 10084
rect 11572 10112 11578 10124
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11572 10084 11897 10112
rect 11572 10072 11578 10084
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 16592 10121 16620 10220
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 18196 10220 18245 10248
rect 18196 10208 18202 10220
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 18233 10211 18291 10217
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12492 10084 13277 10112
rect 12492 10072 12498 10084
rect 13265 10081 13277 10084
rect 13311 10112 13323 10115
rect 13909 10115 13967 10121
rect 13909 10112 13921 10115
rect 13311 10084 13921 10112
rect 13311 10081 13323 10084
rect 13265 10075 13323 10081
rect 13909 10081 13921 10084
rect 13955 10112 13967 10115
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 13955 10084 14105 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 16577 10115 16635 10121
rect 16577 10081 16589 10115
rect 16623 10081 16635 10115
rect 16577 10075 16635 10081
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18104 10084 18521 10112
rect 18104 10072 18110 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 18509 10075 18567 10081
rect 18690 10072 18696 10124
rect 18748 10072 18754 10124
rect 20438 10072 20444 10124
rect 20496 10072 20502 10124
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8202 10044 8208 10056
rect 8067 10016 8208 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 4971 9948 5120 9976
rect 5169 9979 5227 9985
rect 4971 9945 4983 9948
rect 4925 9939 4983 9945
rect 5169 9945 5181 9979
rect 5215 9976 5227 9979
rect 5258 9976 5264 9988
rect 5215 9948 5264 9976
rect 5215 9945 5227 9948
rect 5169 9939 5227 9945
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 5353 9979 5411 9985
rect 5353 9945 5365 9979
rect 5399 9976 5411 9979
rect 6086 9976 6092 9988
rect 5399 9948 6092 9976
rect 5399 9945 5411 9948
rect 5353 9939 5411 9945
rect 6086 9936 6092 9948
rect 6144 9936 6150 9988
rect 6454 9936 6460 9988
rect 6512 9976 6518 9988
rect 6512 9948 6578 9976
rect 6512 9936 6518 9948
rect 7742 9936 7748 9988
rect 7800 9976 7806 9988
rect 8036 9976 8064 10007
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9214 10004 9220 10056
rect 9272 10004 9278 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9490 10044 9496 10056
rect 9447 10016 9496 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10318 10044 10324 10056
rect 9732 10016 10324 10044
rect 9732 10004 9738 10016
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 12158 10004 12164 10056
rect 12216 10004 12222 10056
rect 16844 10047 16902 10053
rect 16844 10013 16856 10047
rect 16890 10044 16902 10047
rect 18322 10044 18328 10056
rect 16890 10016 18328 10044
rect 16890 10013 16902 10016
rect 16844 10007 16902 10013
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 20165 10047 20223 10053
rect 20165 10013 20177 10047
rect 20211 10013 20223 10047
rect 20165 10007 20223 10013
rect 7800 9948 8064 9976
rect 8573 9979 8631 9985
rect 7800 9936 7806 9948
rect 8573 9945 8585 9979
rect 8619 9945 8631 9979
rect 8573 9939 8631 9945
rect 8757 9979 8815 9985
rect 8757 9945 8769 9979
rect 8803 9976 8815 9979
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8803 9948 8953 9976
rect 8803 9945 8815 9948
rect 8757 9939 8815 9945
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 11178 9948 11284 9976
rect 8941 9939 8999 9945
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9877 3663 9911
rect 3605 9871 3663 9877
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4157 9911 4215 9917
rect 4157 9908 4169 9911
rect 4120 9880 4169 9908
rect 4120 9868 4126 9880
rect 4157 9877 4169 9880
rect 4203 9908 4215 9911
rect 5074 9908 5080 9920
rect 4203 9880 5080 9908
rect 4203 9877 4215 9880
rect 4157 9871 4215 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 8588 9908 8616 9939
rect 9306 9908 9312 9920
rect 8588 9880 9312 9908
rect 9306 9868 9312 9880
rect 9364 9908 9370 9920
rect 10042 9908 10048 9920
rect 9364 9880 10048 9908
rect 9364 9868 9370 9880
rect 10042 9868 10048 9880
rect 10100 9908 10106 9920
rect 10137 9911 10195 9917
rect 10137 9908 10149 9911
rect 10100 9880 10149 9908
rect 10100 9868 10106 9880
rect 10137 9877 10149 9880
rect 10183 9877 10195 9911
rect 11256 9908 11284 9948
rect 11606 9936 11612 9988
rect 11664 9936 11670 9988
rect 12176 9908 12204 10004
rect 14366 9985 14372 9988
rect 14360 9976 14372 9985
rect 14327 9948 14372 9976
rect 14360 9939 14372 9948
rect 14366 9936 14372 9939
rect 14424 9936 14430 9988
rect 18785 9979 18843 9985
rect 18785 9976 18797 9979
rect 17972 9948 18797 9976
rect 17972 9920 18000 9948
rect 18785 9945 18797 9948
rect 18831 9945 18843 9979
rect 18785 9939 18843 9945
rect 18874 9936 18880 9988
rect 18932 9976 18938 9988
rect 20180 9976 20208 10007
rect 18932 9948 20208 9976
rect 18932 9936 18938 9948
rect 11256 9880 12204 9908
rect 10137 9871 10195 9877
rect 17954 9868 17960 9920
rect 18012 9868 18018 9920
rect 1104 9818 20792 9840
rect 1104 9766 7214 9818
rect 7266 9766 7278 9818
rect 7330 9766 7342 9818
rect 7394 9766 7406 9818
rect 7458 9766 7470 9818
rect 7522 9766 13214 9818
rect 13266 9766 13278 9818
rect 13330 9766 13342 9818
rect 13394 9766 13406 9818
rect 13458 9766 13470 9818
rect 13522 9766 19214 9818
rect 19266 9766 19278 9818
rect 19330 9766 19342 9818
rect 19394 9766 19406 9818
rect 19458 9766 19470 9818
rect 19522 9766 20792 9818
rect 1104 9744 20792 9766
rect 2498 9664 2504 9716
rect 2556 9664 2562 9716
rect 6457 9707 6515 9713
rect 6457 9673 6469 9707
rect 6503 9704 6515 9707
rect 6546 9704 6552 9716
rect 6503 9676 6552 9704
rect 6503 9673 6515 9676
rect 6457 9667 6515 9673
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 7742 9664 7748 9716
rect 7800 9664 7806 9716
rect 8113 9707 8171 9713
rect 8113 9704 8125 9707
rect 7852 9676 8125 9704
rect 2516 9636 2544 9664
rect 3786 9636 3792 9648
rect 2516 9608 3792 9636
rect 3786 9596 3792 9608
rect 3844 9636 3850 9648
rect 5534 9636 5540 9648
rect 3844 9608 5540 9636
rect 3844 9596 3850 9608
rect 5534 9596 5540 9608
rect 5592 9636 5598 9648
rect 6181 9639 6239 9645
rect 6181 9636 6193 9639
rect 5592 9608 6193 9636
rect 5592 9596 5598 9608
rect 6181 9605 6193 9608
rect 6227 9636 6239 9639
rect 6270 9636 6276 9648
rect 6227 9608 6276 9636
rect 6227 9605 6239 9608
rect 6181 9599 6239 9605
rect 6270 9596 6276 9608
rect 6328 9636 6334 9648
rect 7760 9636 7788 9664
rect 6328 9608 7788 9636
rect 6328 9596 6334 9608
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9568 1639 9571
rect 1670 9568 1676 9580
rect 1627 9540 1676 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6144 9540 6316 9568
rect 6144 9528 6150 9540
rect 6288 9500 6316 9540
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6472 9540 6561 9568
rect 6472 9500 6500 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6788 9540 6868 9568
rect 6788 9528 6794 9540
rect 6288 9472 6500 9500
rect 5074 9392 5080 9444
rect 5132 9432 5138 9444
rect 6840 9432 6868 9540
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 7852 9568 7880 9676
rect 8113 9673 8125 9676
rect 8159 9673 8171 9707
rect 9766 9704 9772 9716
rect 8113 9667 8171 9673
rect 9232 9676 9772 9704
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 9232 9636 9260 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 10318 9664 10324 9716
rect 10376 9664 10382 9716
rect 15010 9664 15016 9716
rect 15068 9704 15074 9716
rect 15473 9707 15531 9713
rect 15473 9704 15485 9707
rect 15068 9676 15485 9704
rect 15068 9664 15074 9676
rect 15473 9673 15485 9676
rect 15519 9673 15531 9707
rect 15473 9667 15531 9673
rect 17497 9707 17555 9713
rect 17497 9673 17509 9707
rect 17543 9704 17555 9707
rect 18414 9704 18420 9716
rect 17543 9676 18420 9704
rect 17543 9673 17555 9676
rect 17497 9667 17555 9673
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 8260 9608 9260 9636
rect 8260 9596 8266 9608
rect 7800 9540 7880 9568
rect 7800 9528 7806 9540
rect 7926 9528 7932 9580
rect 7984 9528 7990 9580
rect 8021 9574 8079 9577
rect 8110 9574 8116 9580
rect 8021 9571 8116 9574
rect 8021 9537 8033 9571
rect 8067 9546 8116 9571
rect 8067 9537 8079 9546
rect 8021 9531 8079 9537
rect 8036 9432 8064 9531
rect 8110 9528 8116 9546
rect 8168 9528 8174 9580
rect 8588 9577 8616 9608
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 17773 9639 17831 9645
rect 17773 9636 17785 9639
rect 14424 9608 17785 9636
rect 14424 9596 14430 9608
rect 17773 9605 17785 9608
rect 17819 9636 17831 9639
rect 18874 9636 18880 9648
rect 17819 9608 18880 9636
rect 17819 9605 17831 9608
rect 17773 9599 17831 9605
rect 18874 9596 18880 9608
rect 18932 9596 18938 9648
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9568 8447 9571
rect 8573 9571 8631 9577
rect 8435 9540 8524 9568
rect 8435 9537 8447 9540
rect 8389 9531 8447 9537
rect 8496 9512 8524 9540
rect 8573 9537 8585 9571
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 14182 9568 14188 9580
rect 10008 9540 14188 9568
rect 10008 9528 10014 9540
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 17681 9571 17739 9577
rect 17681 9537 17693 9571
rect 17727 9568 17739 9571
rect 17954 9568 17960 9580
rect 17727 9540 17960 9568
rect 17727 9537 17739 9540
rect 17681 9531 17739 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18141 9571 18199 9577
rect 18141 9537 18153 9571
rect 18187 9568 18199 9571
rect 18322 9568 18328 9580
rect 18187 9540 18328 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18322 9528 18328 9540
rect 18380 9528 18386 9580
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9568 18475 9571
rect 19714 9571 19772 9577
rect 19714 9568 19726 9571
rect 18463 9540 19726 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 18892 9512 18920 9540
rect 19714 9537 19726 9540
rect 19760 9537 19772 9571
rect 19714 9531 19772 9537
rect 19981 9571 20039 9577
rect 19981 9537 19993 9571
rect 20027 9568 20039 9571
rect 20070 9568 20076 9580
rect 20027 9540 20076 9568
rect 20027 9537 20039 9540
rect 19981 9531 20039 9537
rect 20070 9528 20076 9540
rect 20128 9528 20134 9580
rect 8294 9509 8300 9512
rect 8251 9503 8300 9509
rect 8251 9469 8263 9503
rect 8297 9469 8300 9503
rect 8251 9463 8300 9469
rect 8294 9460 8300 9463
rect 8352 9460 8358 9512
rect 8478 9460 8484 9512
rect 8536 9460 8542 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 8588 9472 8861 9500
rect 8588 9432 8616 9472
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18288 9472 18644 9500
rect 18288 9460 18294 9472
rect 18616 9441 18644 9472
rect 18874 9460 18880 9512
rect 18932 9460 18938 9512
rect 5132 9404 8064 9432
rect 8496 9404 8616 9432
rect 17589 9435 17647 9441
rect 5132 9392 5138 9404
rect 2222 9324 2228 9376
rect 2280 9324 2286 9376
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 6638 9364 6644 9376
rect 4856 9336 6644 9364
rect 4856 9324 4862 9336
rect 6638 9324 6644 9336
rect 6696 9364 6702 9376
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 6696 9336 6745 9364
rect 6696 9324 6702 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 8389 9367 8447 9373
rect 8389 9333 8401 9367
rect 8435 9364 8447 9367
rect 8496 9364 8524 9404
rect 17589 9401 17601 9435
rect 17635 9432 17647 9435
rect 17957 9435 18015 9441
rect 17957 9432 17969 9435
rect 17635 9404 17969 9432
rect 17635 9401 17647 9404
rect 17589 9395 17647 9401
rect 17957 9401 17969 9404
rect 18003 9401 18015 9435
rect 17957 9395 18015 9401
rect 18601 9435 18659 9441
rect 18601 9401 18613 9435
rect 18647 9432 18659 9435
rect 18782 9432 18788 9444
rect 18647 9404 18788 9432
rect 18647 9401 18659 9404
rect 18601 9395 18659 9401
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 8435 9336 8524 9364
rect 8435 9333 8447 9336
rect 8389 9327 8447 9333
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 9858 9364 9864 9376
rect 8628 9336 9864 9364
rect 8628 9324 8634 9336
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 18417 9367 18475 9373
rect 18417 9333 18429 9367
rect 18463 9364 18475 9367
rect 18506 9364 18512 9376
rect 18463 9336 18512 9364
rect 18463 9333 18475 9336
rect 18417 9327 18475 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 1104 9274 20792 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 10214 9274
rect 10266 9222 10278 9274
rect 10330 9222 10342 9274
rect 10394 9222 10406 9274
rect 10458 9222 10470 9274
rect 10522 9222 16214 9274
rect 16266 9222 16278 9274
rect 16330 9222 16342 9274
rect 16394 9222 16406 9274
rect 16458 9222 16470 9274
rect 16522 9222 20792 9274
rect 1104 9200 20792 9222
rect 2222 9120 2228 9172
rect 2280 9120 2286 9172
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 6178 9160 6184 9172
rect 3384 9132 6184 9160
rect 3384 9120 3390 9132
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6270 9120 6276 9172
rect 6328 9120 6334 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8757 9163 8815 9169
rect 8757 9160 8769 9163
rect 8352 9132 8769 9160
rect 8352 9120 8358 9132
rect 8757 9129 8769 9132
rect 8803 9129 8815 9163
rect 8757 9123 8815 9129
rect 17402 9120 17408 9172
rect 17460 9120 17466 9172
rect 17773 9163 17831 9169
rect 17773 9129 17785 9163
rect 17819 9160 17831 9163
rect 17954 9160 17960 9172
rect 17819 9132 17960 9160
rect 17819 9129 17831 9132
rect 17773 9123 17831 9129
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18690 9120 18696 9172
rect 18748 9160 18754 9172
rect 19061 9163 19119 9169
rect 19061 9160 19073 9163
rect 18748 9132 19073 9160
rect 18748 9120 18754 9132
rect 19061 9129 19073 9132
rect 19107 9129 19119 9163
rect 19061 9123 19119 9129
rect 20070 9120 20076 9172
rect 20128 9120 20134 9172
rect 2240 8956 2268 9120
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 8478 9092 8484 9104
rect 6972 9064 8484 9092
rect 6972 9052 6978 9064
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 17862 9092 17868 9104
rect 17144 9064 17868 9092
rect 4430 8984 4436 9036
rect 4488 9024 4494 9036
rect 5074 9024 5080 9036
rect 4488 8996 5080 9024
rect 4488 8984 4494 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5258 8984 5264 9036
rect 5316 8984 5322 9036
rect 7116 8996 7604 9024
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 2240 8928 2329 8956
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8956 5043 8959
rect 5276 8956 5304 8984
rect 5031 8928 5304 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 7116 8965 7144 8996
rect 7576 8968 7604 8996
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 17144 9033 17172 9064
rect 17862 9052 17868 9064
rect 17920 9092 17926 9104
rect 18325 9095 18383 9101
rect 18325 9092 18337 9095
rect 17920 9064 18337 9092
rect 17920 9052 17926 9064
rect 18325 9061 18337 9064
rect 18371 9092 18383 9095
rect 18966 9092 18972 9104
rect 18371 9064 18972 9092
rect 18371 9061 18383 9064
rect 18325 9055 18383 9061
rect 18966 9052 18972 9064
rect 19024 9092 19030 9104
rect 20088 9092 20116 9120
rect 19024 9064 20116 9092
rect 19024 9052 19030 9064
rect 17129 9027 17187 9033
rect 7800 8996 8800 9024
rect 7800 8984 7806 8996
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 4893 8891 4951 8897
rect 4893 8857 4905 8891
rect 4939 8888 4951 8891
rect 6380 8888 6408 8916
rect 4939 8860 6408 8888
rect 4939 8857 4951 8860
rect 4893 8851 4951 8857
rect 5000 8832 5028 8860
rect 6730 8848 6736 8900
rect 6788 8888 6794 8900
rect 7392 8888 7420 8919
rect 7558 8916 7564 8968
rect 7616 8916 7622 8968
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7668 8928 7849 8956
rect 6788 8860 7420 8888
rect 6788 8848 6794 8860
rect 7668 8832 7696 8928
rect 7837 8925 7849 8928
rect 7883 8956 7895 8959
rect 7926 8956 7932 8968
rect 7883 8928 7932 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 7926 8916 7932 8928
rect 7984 8956 7990 8968
rect 8772 8965 8800 8996
rect 17129 8993 17141 9027
rect 17175 8993 17187 9027
rect 17129 8987 17187 8993
rect 18506 8984 18512 9036
rect 18564 9024 18570 9036
rect 18564 8996 18736 9024
rect 18564 8984 18570 8996
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 7984 8928 8493 8956
rect 7984 8916 7990 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9674 8956 9680 8968
rect 8803 8928 9680 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 10597 8959 10655 8965
rect 10597 8925 10609 8959
rect 10643 8925 10655 8959
rect 10597 8919 10655 8925
rect 13909 8959 13967 8965
rect 13909 8925 13921 8959
rect 13955 8956 13967 8959
rect 14090 8956 14096 8968
rect 13955 8928 14096 8956
rect 13955 8925 13967 8928
rect 13909 8919 13967 8925
rect 1670 8780 1676 8832
rect 1728 8780 1734 8832
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4396 8792 4537 8820
rect 4396 8780 4402 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 4982 8780 4988 8832
rect 5040 8780 5046 8832
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 7006 8820 7012 8832
rect 6963 8792 7012 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 7006 8780 7012 8792
rect 7064 8780 7070 8832
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 7156 8792 7297 8820
rect 7156 8780 7162 8792
rect 7285 8789 7297 8792
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 7650 8780 7656 8832
rect 7708 8780 7714 8832
rect 7742 8780 7748 8832
rect 7800 8780 7806 8832
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8570 8820 8576 8832
rect 8168 8792 8576 8820
rect 8168 8780 8174 8792
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 10612 8820 10640 8919
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 14366 8965 14372 8968
rect 14360 8919 14372 8965
rect 14366 8916 14372 8919
rect 14424 8916 14430 8968
rect 17586 8916 17592 8968
rect 17644 8916 17650 8968
rect 18708 8965 18736 8996
rect 17773 8959 17831 8965
rect 17773 8925 17785 8959
rect 17819 8925 17831 8959
rect 17773 8919 17831 8925
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 18693 8919 18751 8925
rect 10778 8848 10784 8900
rect 10836 8888 10842 8900
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 10836 8860 10885 8888
rect 10836 8848 10842 8860
rect 10873 8857 10885 8860
rect 10919 8857 10931 8891
rect 13722 8888 13728 8900
rect 12098 8860 13728 8888
rect 10873 8851 10931 8857
rect 13722 8848 13728 8860
rect 13780 8848 13786 8900
rect 16850 8848 16856 8900
rect 16908 8897 16914 8900
rect 16908 8851 16920 8897
rect 17788 8888 17816 8919
rect 17788 8860 18460 8888
rect 16908 8848 16914 8851
rect 11054 8820 11060 8832
rect 10612 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 12345 8823 12403 8829
rect 12345 8820 12357 8823
rect 12216 8792 12357 8820
rect 12216 8780 12222 8792
rect 12345 8789 12357 8792
rect 12391 8789 12403 8823
rect 12345 8783 12403 8789
rect 15470 8780 15476 8832
rect 15528 8780 15534 8832
rect 15746 8780 15752 8832
rect 15804 8780 15810 8832
rect 18432 8820 18460 8860
rect 18506 8848 18512 8900
rect 18564 8848 18570 8900
rect 20346 8888 20352 8900
rect 18708 8860 20352 8888
rect 18708 8820 18736 8860
rect 20346 8848 20352 8860
rect 20404 8848 20410 8900
rect 18432 8792 18736 8820
rect 18782 8780 18788 8832
rect 18840 8780 18846 8832
rect 18874 8780 18880 8832
rect 18932 8780 18938 8832
rect 1104 8730 20792 8752
rect 1104 8678 7214 8730
rect 7266 8678 7278 8730
rect 7330 8678 7342 8730
rect 7394 8678 7406 8730
rect 7458 8678 7470 8730
rect 7522 8678 13214 8730
rect 13266 8678 13278 8730
rect 13330 8678 13342 8730
rect 13394 8678 13406 8730
rect 13458 8678 13470 8730
rect 13522 8678 19214 8730
rect 19266 8678 19278 8730
rect 19330 8678 19342 8730
rect 19394 8678 19406 8730
rect 19458 8678 19470 8730
rect 19522 8678 20792 8730
rect 1104 8656 20792 8678
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8616 3755 8619
rect 3786 8616 3792 8628
rect 3743 8588 3792 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 4338 8616 4344 8628
rect 4172 8588 4344 8616
rect 4172 8557 4200 8588
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4430 8576 4436 8628
rect 4488 8576 4494 8628
rect 4798 8616 4804 8628
rect 4540 8588 4804 8616
rect 4157 8551 4215 8557
rect 4157 8517 4169 8551
rect 4203 8517 4215 8551
rect 4157 8511 4215 8517
rect 4249 8551 4307 8557
rect 4249 8517 4261 8551
rect 4295 8548 4307 8551
rect 4448 8548 4476 8576
rect 4295 8520 4476 8548
rect 4295 8517 4307 8520
rect 4249 8511 4307 8517
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4367 8483 4425 8489
rect 4367 8449 4379 8483
rect 4413 8480 4425 8483
rect 4540 8480 4568 8588
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 5258 8616 5264 8628
rect 5092 8588 5264 8616
rect 4982 8548 4988 8560
rect 4632 8520 4988 8548
rect 4632 8489 4660 8520
rect 4982 8508 4988 8520
rect 5040 8508 5046 8560
rect 4413 8452 4568 8480
rect 4617 8483 4675 8489
rect 4413 8449 4425 8452
rect 4367 8443 4425 8449
rect 4617 8449 4629 8483
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 4080 8344 4108 8443
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 4893 8483 4951 8489
rect 4764 8452 4844 8480
rect 4764 8440 4770 8452
rect 4154 8372 4160 8424
rect 4212 8412 4218 8424
rect 4525 8415 4583 8421
rect 4525 8412 4537 8415
rect 4212 8384 4537 8412
rect 4212 8372 4218 8384
rect 4525 8381 4537 8384
rect 4571 8412 4583 8415
rect 4816 8412 4844 8452
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 5092 8480 5120 8588
rect 5258 8576 5264 8588
rect 5316 8616 5322 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 5316 8588 5365 8616
rect 5316 8576 5322 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 5353 8579 5411 8585
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5718 8616 5724 8628
rect 5675 8588 5724 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 10505 8619 10563 8625
rect 6236 8588 10456 8616
rect 6236 8576 6242 8588
rect 5184 8520 5856 8548
rect 5184 8489 5212 8520
rect 5828 8489 5856 8520
rect 7466 8508 7472 8560
rect 7524 8508 7530 8560
rect 9306 8508 9312 8560
rect 9364 8508 9370 8560
rect 4939 8452 5120 8480
rect 5169 8483 5227 8489
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 5169 8449 5181 8483
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8480 6147 8483
rect 6178 8480 6184 8492
rect 6135 8452 6184 8480
rect 6135 8449 6147 8452
rect 6089 8443 6147 8449
rect 5184 8412 5212 8443
rect 4571 8384 5212 8412
rect 5276 8412 5304 8443
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 10428 8489 10456 8588
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 10778 8616 10784 8628
rect 10551 8588 10784 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11054 8576 11060 8628
rect 11112 8576 11118 8628
rect 11238 8576 11244 8628
rect 11296 8625 11302 8628
rect 11296 8616 11307 8625
rect 12434 8616 12440 8628
rect 11296 8588 11341 8616
rect 11296 8579 11307 8588
rect 11296 8576 11302 8579
rect 12406 8576 12440 8616
rect 12492 8576 12498 8628
rect 16317 8619 16375 8625
rect 16317 8616 16329 8619
rect 15488 8588 16329 8616
rect 10873 8551 10931 8557
rect 10873 8517 10885 8551
rect 10919 8548 10931 8551
rect 11072 8548 11100 8576
rect 12406 8548 12434 8576
rect 15488 8560 15516 8588
rect 16317 8585 16329 8588
rect 16363 8616 16375 8619
rect 16485 8619 16543 8625
rect 16363 8588 16436 8616
rect 16363 8585 16375 8588
rect 16317 8579 16375 8585
rect 10919 8520 11652 8548
rect 10919 8517 10931 8520
rect 10873 8511 10931 8517
rect 11624 8492 11652 8520
rect 11992 8520 12434 8548
rect 13832 8520 14582 8548
rect 6457 8483 6515 8489
rect 6457 8480 6469 8483
rect 6328 8452 6469 8480
rect 6328 8440 6334 8452
rect 6457 8449 6469 8452
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10413 8443 10471 8449
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 10597 8443 10655 8449
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8480 10747 8483
rect 10778 8480 10784 8492
rect 10735 8452 10784 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 5276 8384 5396 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 5368 8344 5396 8384
rect 5902 8372 5908 8424
rect 5960 8372 5966 8424
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8412 6791 8415
rect 7282 8412 7288 8424
rect 6779 8384 7288 8412
rect 6779 8381 6791 8384
rect 6733 8375 6791 8381
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8536 8384 8953 8412
rect 8536 8372 8542 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 4080 8316 4844 8344
rect 5368 8316 5672 8344
rect 2406 8236 2412 8288
rect 2464 8236 2470 8288
rect 3878 8236 3884 8288
rect 3936 8236 3942 8288
rect 4816 8285 4844 8316
rect 4801 8279 4859 8285
rect 4801 8245 4813 8279
rect 4847 8276 4859 8279
rect 5166 8276 5172 8288
rect 4847 8248 5172 8276
rect 4847 8245 4859 8248
rect 4801 8239 4859 8245
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5534 8236 5540 8288
rect 5592 8236 5598 8288
rect 5644 8276 5672 8316
rect 7742 8304 7748 8356
rect 7800 8304 7806 8356
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8389 8347 8447 8353
rect 8389 8344 8401 8347
rect 8352 8316 8401 8344
rect 8352 8304 8358 8316
rect 8389 8313 8401 8316
rect 8435 8313 8447 8347
rect 8389 8307 8447 8313
rect 9674 8304 9680 8356
rect 9732 8304 9738 8356
rect 10428 8344 10456 8443
rect 10612 8412 10640 8443
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 11109 8483 11167 8489
rect 11109 8449 11121 8483
rect 11155 8480 11167 8483
rect 11155 8452 11560 8480
rect 11155 8449 11167 8452
rect 11109 8443 11167 8449
rect 10980 8412 11008 8443
rect 10612 8384 11008 8412
rect 11532 8412 11560 8452
rect 11606 8440 11612 8492
rect 11664 8440 11670 8492
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 11992 8421 12020 8520
rect 13722 8480 13728 8492
rect 13386 8452 13728 8480
rect 13722 8440 13728 8452
rect 13780 8480 13786 8492
rect 13832 8480 13860 8520
rect 15470 8508 15476 8560
rect 15528 8508 15534 8560
rect 15746 8508 15752 8560
rect 15804 8548 15810 8560
rect 16117 8551 16175 8557
rect 16117 8548 16129 8551
rect 15804 8520 16129 8548
rect 15804 8508 15810 8520
rect 16117 8517 16129 8520
rect 16163 8517 16175 8551
rect 16117 8511 16175 8517
rect 13780 8452 13860 8480
rect 13780 8440 13786 8452
rect 11977 8415 12035 8421
rect 11977 8412 11989 8415
rect 11532 8384 11989 8412
rect 10980 8344 11008 8384
rect 11977 8381 11989 8384
rect 12023 8381 12035 8415
rect 11977 8375 12035 8381
rect 12084 8384 13768 8412
rect 12084 8344 12112 8384
rect 10428 8316 10916 8344
rect 10980 8316 12112 8344
rect 13740 8344 13768 8384
rect 13814 8372 13820 8424
rect 13872 8372 13878 8424
rect 15565 8415 15623 8421
rect 15565 8412 15577 8415
rect 13924 8384 15577 8412
rect 13924 8344 13952 8384
rect 15565 8381 15577 8384
rect 15611 8381 15623 8415
rect 16132 8412 16160 8511
rect 16408 8480 16436 8588
rect 16485 8585 16497 8619
rect 16531 8585 16543 8619
rect 16485 8579 16543 8585
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 17586 8616 17592 8628
rect 17083 8588 17592 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 16500 8548 16528 8579
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 17221 8551 17279 8557
rect 17221 8548 17233 8551
rect 16500 8520 17233 8548
rect 17221 8517 17233 8520
rect 17267 8517 17279 8551
rect 17221 8511 17279 8517
rect 17437 8551 17495 8557
rect 17437 8517 17449 8551
rect 17483 8548 17495 8551
rect 19242 8548 19248 8560
rect 17483 8520 19248 8548
rect 17483 8517 17495 8520
rect 17437 8511 17495 8517
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 16408 8452 16681 8480
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 17862 8440 17868 8492
rect 17920 8440 17926 8492
rect 18138 8489 18144 8492
rect 18132 8480 18144 8489
rect 18099 8452 18144 8480
rect 18132 8443 18144 8452
rect 18138 8440 18144 8443
rect 18196 8440 18202 8492
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 16132 8384 16773 8412
rect 15565 8375 15623 8381
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 16761 8375 16819 8381
rect 13740 8316 13952 8344
rect 17589 8347 17647 8353
rect 5810 8276 5816 8288
rect 5644 8248 5816 8276
rect 5810 8236 5816 8248
rect 5868 8236 5874 8288
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 7760 8276 7788 8304
rect 7248 8248 7788 8276
rect 7248 8236 7254 8248
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7892 8248 8217 8276
rect 7892 8236 7898 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8205 8239 8263 8245
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 9125 8279 9183 8285
rect 9125 8276 9137 8279
rect 8996 8248 9137 8276
rect 8996 8236 9002 8248
rect 9125 8245 9137 8248
rect 9171 8245 9183 8279
rect 9125 8239 9183 8245
rect 9309 8279 9367 8285
rect 9309 8245 9321 8279
rect 9355 8276 9367 8279
rect 9582 8276 9588 8288
rect 9355 8248 9588 8276
rect 9355 8245 9367 8248
rect 9309 8239 9367 8245
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 10888 8276 10916 8316
rect 17589 8313 17601 8347
rect 17635 8344 17647 8347
rect 18892 8344 18920 8440
rect 19245 8347 19303 8353
rect 19245 8344 19257 8347
rect 17635 8316 17908 8344
rect 18892 8316 19257 8344
rect 17635 8313 17647 8316
rect 17589 8307 17647 8313
rect 11330 8276 11336 8288
rect 10888 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11885 8279 11943 8285
rect 11885 8245 11897 8279
rect 11931 8276 11943 8279
rect 12234 8279 12292 8285
rect 12234 8276 12246 8279
rect 11931 8248 12246 8276
rect 11931 8245 11943 8248
rect 11885 8239 11943 8245
rect 12234 8245 12246 8248
rect 12280 8245 12292 8279
rect 12234 8239 12292 8245
rect 13725 8279 13783 8285
rect 13725 8245 13737 8279
rect 13771 8276 13783 8279
rect 14074 8279 14132 8285
rect 14074 8276 14086 8279
rect 13771 8248 14086 8276
rect 13771 8245 13783 8248
rect 13725 8239 13783 8245
rect 14074 8245 14086 8248
rect 14120 8245 14132 8279
rect 14074 8239 14132 8245
rect 16301 8279 16359 8285
rect 16301 8245 16313 8279
rect 16347 8276 16359 8279
rect 16850 8276 16856 8288
rect 16347 8248 16856 8276
rect 16347 8245 16359 8248
rect 16301 8239 16359 8245
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 17402 8236 17408 8288
rect 17460 8236 17466 8288
rect 17880 8276 17908 8316
rect 19245 8313 19257 8316
rect 19291 8313 19303 8347
rect 19245 8307 19303 8313
rect 18046 8276 18052 8288
rect 17880 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 1104 8186 20792 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 10214 8186
rect 10266 8134 10278 8186
rect 10330 8134 10342 8186
rect 10394 8134 10406 8186
rect 10458 8134 10470 8186
rect 10522 8134 16214 8186
rect 16266 8134 16278 8186
rect 16330 8134 16342 8186
rect 16394 8134 16406 8186
rect 16458 8134 16470 8186
rect 16522 8134 20792 8186
rect 1104 8112 20792 8134
rect 2120 8075 2178 8081
rect 2120 8041 2132 8075
rect 2166 8072 2178 8075
rect 3878 8072 3884 8084
rect 2166 8044 3884 8072
rect 2166 8041 2178 8044
rect 2120 8035 2178 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 5408 8044 5549 8072
rect 5408 8032 5414 8044
rect 5537 8041 5549 8044
rect 5583 8072 5595 8075
rect 5810 8072 5816 8084
rect 5583 8044 5816 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6730 8072 6736 8084
rect 5920 8044 6736 8072
rect 5920 8004 5948 8044
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7282 8032 7288 8084
rect 7340 8032 7346 8084
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7708 8044 7757 8072
rect 7708 8032 7714 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 7834 8032 7840 8084
rect 7892 8032 7898 8084
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 11517 8075 11575 8081
rect 8260 8044 10732 8072
rect 8260 8032 8266 8044
rect 3620 7976 3924 8004
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 2222 7936 2228 7948
rect 1903 7908 2228 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 2222 7896 2228 7908
rect 2280 7936 2286 7948
rect 2498 7936 2504 7948
rect 2280 7908 2504 7936
rect 2280 7896 2286 7908
rect 2498 7896 2504 7908
rect 2556 7936 2562 7948
rect 3142 7936 3148 7948
rect 2556 7908 3148 7936
rect 2556 7896 2562 7908
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 3620 7868 3648 7976
rect 3789 7939 3847 7945
rect 3789 7905 3801 7939
rect 3835 7905 3847 7939
rect 3896 7936 3924 7976
rect 5644 7976 5948 8004
rect 4798 7936 4804 7948
rect 3896 7908 4804 7936
rect 3789 7899 3847 7905
rect 3266 7840 3648 7868
rect 3694 7800 3700 7812
rect 3528 7772 3700 7800
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 3528 7732 3556 7772
rect 3694 7760 3700 7772
rect 3752 7800 3758 7812
rect 3804 7800 3832 7899
rect 4798 7896 4804 7908
rect 4856 7896 4862 7948
rect 5534 7896 5540 7948
rect 5592 7936 5598 7948
rect 5644 7936 5672 7976
rect 6178 7964 6184 8016
rect 6236 8004 6242 8016
rect 7576 8004 7604 8032
rect 7852 8004 7880 8032
rect 6236 7976 7880 8004
rect 6236 7964 6242 7976
rect 6656 7945 6684 7976
rect 6365 7939 6423 7945
rect 6365 7936 6377 7939
rect 5592 7908 5672 7936
rect 5592 7896 5598 7908
rect 5644 7877 5672 7908
rect 5828 7908 6377 7936
rect 5828 7877 5856 7908
rect 6365 7905 6377 7908
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 6730 7896 6736 7948
rect 6788 7936 6794 7948
rect 6788 7908 7512 7936
rect 6788 7896 6794 7908
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 5994 7828 6000 7880
rect 6052 7828 6058 7880
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 6144 7840 6285 7868
rect 6144 7828 6150 7840
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 3752 7772 3832 7800
rect 3752 7760 3758 7772
rect 4062 7760 4068 7812
rect 4120 7760 4126 7812
rect 4798 7760 4804 7812
rect 4856 7760 4862 7812
rect 5902 7760 5908 7812
rect 5960 7800 5966 7812
rect 6472 7800 6500 7831
rect 7006 7828 7012 7880
rect 7064 7828 7070 7880
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7868 7159 7871
rect 7190 7868 7196 7880
rect 7147 7840 7196 7868
rect 7147 7837 7159 7840
rect 7101 7831 7159 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7484 7862 7512 7908
rect 7558 7896 7564 7948
rect 7616 7936 7622 7948
rect 8665 7939 8723 7945
rect 8665 7936 8677 7939
rect 7616 7908 8677 7936
rect 7616 7896 7622 7908
rect 8665 7905 8677 7908
rect 8711 7905 8723 7939
rect 8665 7899 8723 7905
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 9674 7936 9680 7948
rect 8987 7908 9680 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10704 7945 10732 8044
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 11698 8072 11704 8084
rect 11563 8044 11704 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 13725 8075 13783 8081
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 13814 8072 13820 8084
rect 13771 8044 13820 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 16117 8075 16175 8081
rect 16117 8041 16129 8075
rect 16163 8072 16175 8075
rect 16850 8072 16856 8084
rect 16163 8044 16856 8072
rect 16163 8041 16175 8044
rect 16117 8035 16175 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 17681 8075 17739 8081
rect 17681 8041 17693 8075
rect 17727 8072 17739 8075
rect 18138 8072 18144 8084
rect 17727 8044 18144 8072
rect 17727 8041 17739 8044
rect 17681 8035 17739 8041
rect 18138 8032 18144 8044
rect 18196 8072 18202 8084
rect 18196 8044 19104 8072
rect 18196 8032 18202 8044
rect 11330 7964 11336 8016
rect 11388 7964 11394 8016
rect 17129 8007 17187 8013
rect 17129 7973 17141 8007
rect 17175 8004 17187 8007
rect 17497 8007 17555 8013
rect 17497 8004 17509 8007
rect 17175 7976 17509 8004
rect 17175 7973 17187 7976
rect 17129 7967 17187 7973
rect 17497 7973 17509 7976
rect 17543 8004 17555 8007
rect 17862 8004 17868 8016
rect 17543 7976 17868 8004
rect 17543 7973 17555 7976
rect 17497 7967 17555 7973
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 19076 8004 19104 8044
rect 19242 8032 19248 8084
rect 19300 8032 19306 8084
rect 20165 8075 20223 8081
rect 20165 8041 20177 8075
rect 20211 8072 20223 8075
rect 20211 8044 20300 8072
rect 20211 8041 20223 8044
rect 20165 8035 20223 8041
rect 19797 8007 19855 8013
rect 19797 8004 19809 8007
rect 19076 7976 19809 8004
rect 19797 7973 19809 7976
rect 19843 8004 19855 8007
rect 19843 7976 20208 8004
rect 19843 7973 19855 7976
rect 19797 7967 19855 7973
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7905 10747 7939
rect 10689 7899 10747 7905
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7936 12127 7939
rect 12158 7936 12164 7948
rect 12115 7908 12164 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 12492 7908 13676 7936
rect 12492 7896 12498 7908
rect 7484 7834 7604 7862
rect 5960 7772 6500 7800
rect 5960 7760 5966 7772
rect 3200 7704 3556 7732
rect 3605 7735 3663 7741
rect 3200 7692 3206 7704
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 3970 7732 3976 7744
rect 3651 7704 3976 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 6178 7692 6184 7744
rect 6236 7692 6242 7744
rect 6472 7732 6500 7772
rect 6638 7760 6644 7812
rect 6696 7800 6702 7812
rect 6779 7803 6837 7809
rect 6779 7800 6791 7803
rect 6696 7772 6791 7800
rect 6696 7760 6702 7772
rect 6779 7769 6791 7772
rect 6825 7769 6837 7803
rect 6779 7763 6837 7769
rect 6914 7760 6920 7812
rect 6972 7760 6978 7812
rect 7377 7803 7435 7809
rect 7377 7769 7389 7803
rect 7423 7769 7435 7803
rect 7377 7763 7435 7769
rect 7006 7732 7012 7744
rect 6472 7704 7012 7732
rect 7006 7692 7012 7704
rect 7064 7732 7070 7744
rect 7392 7732 7420 7763
rect 7064 7704 7420 7732
rect 7576 7741 7604 7834
rect 11790 7828 11796 7880
rect 11848 7828 11854 7880
rect 13648 7877 13676 7908
rect 19518 7896 19524 7948
rect 19576 7936 19582 7948
rect 19702 7936 19708 7948
rect 19576 7908 19708 7936
rect 19576 7896 19582 7908
rect 19702 7896 19708 7908
rect 19760 7936 19766 7948
rect 19981 7939 20039 7945
rect 19981 7936 19993 7939
rect 19760 7908 19993 7936
rect 19760 7896 19766 7908
rect 19981 7905 19993 7908
rect 20027 7905 20039 7939
rect 19981 7899 20039 7905
rect 13633 7871 13691 7877
rect 13633 7837 13645 7871
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 14148 7840 14749 7868
rect 14148 7828 14154 7840
rect 14737 7837 14749 7840
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 15004 7871 15062 7877
rect 15004 7837 15016 7871
rect 15050 7868 15062 7871
rect 15470 7868 15476 7880
rect 15050 7840 15476 7868
rect 15050 7837 15062 7840
rect 15004 7831 15062 7837
rect 7926 7760 7932 7812
rect 7984 7800 7990 7812
rect 8389 7803 8447 7809
rect 8389 7800 8401 7803
rect 7984 7772 8401 7800
rect 7984 7760 7990 7772
rect 8389 7769 8401 7772
rect 8435 7800 8447 7803
rect 8478 7800 8484 7812
rect 8435 7772 8484 7800
rect 8435 7769 8447 7772
rect 8389 7763 8447 7769
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 9398 7760 9404 7812
rect 9456 7760 9462 7812
rect 10413 7803 10471 7809
rect 10413 7769 10425 7803
rect 10459 7769 10471 7803
rect 10413 7763 10471 7769
rect 7576 7735 7645 7741
rect 7576 7704 7599 7735
rect 7064 7692 7070 7704
rect 7587 7701 7599 7704
rect 7633 7701 7645 7735
rect 7587 7695 7645 7701
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 10428 7732 10456 7763
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 13722 7800 13728 7812
rect 11112 7772 12434 7800
rect 13294 7772 13728 7800
rect 11112 7760 11118 7772
rect 9640 7704 10456 7732
rect 12406 7732 12434 7772
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 12406 7704 13553 7732
rect 9640 7692 9646 7704
rect 13541 7701 13553 7704
rect 13587 7701 13599 7735
rect 13541 7695 13599 7701
rect 14645 7735 14703 7741
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 14752 7732 14780 7831
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 19061 7871 19119 7877
rect 19061 7868 19073 7871
rect 19024 7840 19073 7868
rect 19024 7828 19030 7840
rect 19061 7837 19073 7840
rect 19107 7837 19119 7871
rect 19061 7831 19119 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7868 19487 7871
rect 19610 7868 19616 7880
rect 19475 7840 19616 7868
rect 19475 7837 19487 7840
rect 19429 7831 19487 7837
rect 19610 7828 19616 7840
rect 19668 7868 19674 7880
rect 20180 7877 20208 7976
rect 19889 7871 19947 7877
rect 19889 7868 19901 7871
rect 19668 7840 19901 7868
rect 19668 7828 19674 7840
rect 19889 7837 19901 7840
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 18598 7760 18604 7812
rect 18656 7800 18662 7812
rect 18816 7803 18874 7809
rect 18816 7800 18828 7803
rect 18656 7772 18828 7800
rect 18656 7760 18662 7772
rect 18816 7769 18828 7772
rect 18862 7800 18874 7803
rect 18862 7772 19656 7800
rect 18862 7769 18874 7772
rect 18816 7763 18874 7769
rect 15010 7732 15016 7744
rect 14691 7704 15016 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 19518 7692 19524 7744
rect 19576 7692 19582 7744
rect 19628 7741 19656 7772
rect 19613 7735 19671 7741
rect 19613 7701 19625 7735
rect 19659 7732 19671 7735
rect 20272 7732 20300 8044
rect 20346 8032 20352 8084
rect 20404 8032 20410 8084
rect 19659 7704 20300 7732
rect 19659 7701 19671 7704
rect 19613 7695 19671 7701
rect 1104 7642 20792 7664
rect 1104 7590 7214 7642
rect 7266 7590 7278 7642
rect 7330 7590 7342 7642
rect 7394 7590 7406 7642
rect 7458 7590 7470 7642
rect 7522 7590 13214 7642
rect 13266 7590 13278 7642
rect 13330 7590 13342 7642
rect 13394 7590 13406 7642
rect 13458 7590 13470 7642
rect 13522 7590 19214 7642
rect 19266 7590 19278 7642
rect 19330 7590 19342 7642
rect 19394 7590 19406 7642
rect 19458 7590 19470 7642
rect 19522 7590 20792 7642
rect 1104 7568 20792 7590
rect 3694 7488 3700 7540
rect 3752 7488 3758 7540
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4525 7531 4583 7537
rect 4525 7528 4537 7531
rect 4120 7500 4537 7528
rect 4120 7488 4126 7500
rect 4525 7497 4537 7500
rect 4571 7497 4583 7531
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 4525 7491 4583 7497
rect 4816 7500 5733 7528
rect 2406 7420 2412 7472
rect 2464 7420 2470 7472
rect 4816 7460 4844 7500
rect 5721 7497 5733 7500
rect 5767 7528 5779 7531
rect 5994 7528 6000 7540
rect 5767 7500 6000 7528
rect 5767 7497 5779 7500
rect 5721 7491 5779 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 6236 7500 6684 7528
rect 6236 7488 6242 7500
rect 6656 7469 6684 7500
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 8570 7528 8576 7540
rect 6972 7500 8576 7528
rect 6972 7488 6978 7500
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 11609 7531 11667 7537
rect 11609 7497 11621 7531
rect 11655 7528 11667 7531
rect 11790 7528 11796 7540
rect 11655 7500 11796 7528
rect 11655 7497 11667 7500
rect 11609 7491 11667 7497
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 18598 7488 18604 7540
rect 18656 7488 18662 7540
rect 18966 7488 18972 7540
rect 19024 7488 19030 7540
rect 4724 7432 4844 7460
rect 4893 7463 4951 7469
rect 4724 7401 4752 7432
rect 4893 7429 4905 7463
rect 4939 7460 4951 7463
rect 5261 7463 5319 7469
rect 5261 7460 5273 7463
rect 4939 7432 5273 7460
rect 4939 7429 4951 7432
rect 4893 7423 4951 7429
rect 5261 7429 5273 7432
rect 5307 7429 5319 7463
rect 5261 7423 5319 7429
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7429 6699 7463
rect 6641 7423 6699 7429
rect 7098 7420 7104 7472
rect 7156 7420 7162 7472
rect 9582 7460 9588 7472
rect 9232 7432 9588 7460
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 1578 7284 1584 7336
rect 1636 7284 1642 7336
rect 4816 7324 4844 7355
rect 5074 7352 5080 7404
rect 5132 7352 5138 7404
rect 5166 7352 5172 7404
rect 5224 7352 5230 7404
rect 5350 7352 5356 7404
rect 5408 7352 5414 7404
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5368 7324 5396 7352
rect 4816 7296 5396 7324
rect 5460 7324 5488 7355
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5592 7364 5641 7392
rect 5592 7352 5598 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6328 7364 6377 7392
rect 6328 7352 6334 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 8938 7392 8944 7404
rect 8803 7364 8944 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9232 7401 9260 7432
rect 9582 7420 9588 7432
rect 9640 7420 9646 7472
rect 10134 7420 10140 7472
rect 10192 7420 10198 7472
rect 15188 7463 15246 7469
rect 15188 7429 15200 7463
rect 15234 7460 15246 7463
rect 15746 7460 15752 7472
rect 15234 7432 15752 7460
rect 15234 7429 15246 7432
rect 15188 7423 15246 7429
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 18414 7420 18420 7472
rect 18472 7460 18478 7472
rect 18984 7460 19012 7488
rect 18472 7432 20024 7460
rect 18472 7420 18478 7432
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9306 7352 9312 7404
rect 9364 7352 9370 7404
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7392 9551 7395
rect 9674 7392 9680 7404
rect 9539 7364 9680 7392
rect 9539 7361 9551 7364
rect 9493 7355 9551 7361
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7392 11575 7395
rect 11606 7392 11612 7404
rect 11563 7364 11612 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7392 14887 7395
rect 14921 7395 14979 7401
rect 14921 7392 14933 7395
rect 14875 7364 14933 7392
rect 14875 7361 14887 7364
rect 14829 7355 14887 7361
rect 14921 7361 14933 7364
rect 14967 7392 14979 7395
rect 15010 7392 15016 7404
rect 14967 7364 15016 7392
rect 14967 7361 14979 7364
rect 14921 7355 14979 7361
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 19702 7352 19708 7404
rect 19760 7401 19766 7404
rect 19996 7401 20024 7432
rect 19760 7392 19772 7401
rect 19981 7395 20039 7401
rect 19760 7364 19805 7392
rect 19760 7355 19772 7364
rect 19981 7361 19993 7395
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 19760 7352 19766 7355
rect 6086 7324 6092 7336
rect 5460 7296 6092 7324
rect 6086 7284 6092 7296
rect 6144 7324 6150 7336
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 6144 7296 8861 7324
rect 6144 7284 6150 7296
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 5905 7191 5963 7197
rect 5905 7157 5917 7191
rect 5951 7188 5963 7191
rect 6638 7188 6644 7200
rect 5951 7160 6644 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 7064 7160 8125 7188
rect 7064 7148 7070 7160
rect 8113 7157 8125 7160
rect 8159 7157 8171 7191
rect 8113 7151 8171 7157
rect 9398 7148 9404 7200
rect 9456 7188 9462 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 9456 7160 10057 7188
rect 9456 7148 9462 7160
rect 10045 7157 10057 7160
rect 10091 7188 10103 7191
rect 13722 7188 13728 7200
rect 10091 7160 13728 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 16301 7191 16359 7197
rect 16301 7188 16313 7191
rect 16172 7160 16313 7188
rect 16172 7148 16178 7160
rect 16301 7157 16313 7160
rect 16347 7157 16359 7191
rect 16301 7151 16359 7157
rect 1104 7098 20792 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 10214 7098
rect 10266 7046 10278 7098
rect 10330 7046 10342 7098
rect 10394 7046 10406 7098
rect 10458 7046 10470 7098
rect 10522 7046 16214 7098
rect 16266 7046 16278 7098
rect 16330 7046 16342 7098
rect 16394 7046 16406 7098
rect 16458 7046 16470 7098
rect 16522 7046 20792 7098
rect 1104 7024 20792 7046
rect 6270 6944 6276 6996
rect 6328 6944 6334 6996
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 17497 6987 17555 6993
rect 17497 6984 17509 6987
rect 17460 6956 17509 6984
rect 17460 6944 17466 6956
rect 17497 6953 17509 6956
rect 17543 6953 17555 6987
rect 17497 6947 17555 6953
rect 17678 6944 17684 6996
rect 17736 6944 17742 6996
rect 18414 6944 18420 6996
rect 18472 6944 18478 6996
rect 15010 6876 15016 6928
rect 15068 6916 15074 6928
rect 16945 6919 17003 6925
rect 16945 6916 16957 6919
rect 15068 6888 15240 6916
rect 15068 6876 15074 6888
rect 2222 6808 2228 6860
rect 2280 6808 2286 6860
rect 15212 6848 15240 6888
rect 16684 6888 16957 6916
rect 16684 6860 16712 6888
rect 16945 6885 16957 6888
rect 16991 6916 17003 6919
rect 16991 6888 17448 6916
rect 16991 6885 17003 6888
rect 16945 6879 17003 6885
rect 15212 6820 15332 6848
rect 12802 6740 12808 6792
rect 12860 6740 12866 6792
rect 15304 6789 15332 6820
rect 16666 6808 16672 6860
rect 16724 6808 16730 6860
rect 17420 6848 17448 6888
rect 17052 6820 17356 6848
rect 17420 6820 17908 6848
rect 15289 6783 15347 6789
rect 15289 6749 15301 6783
rect 15335 6780 15347 6783
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 15335 6752 15393 6780
rect 15335 6749 15347 6752
rect 15289 6743 15347 6749
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 15648 6783 15706 6789
rect 15648 6749 15660 6783
rect 15694 6780 15706 6783
rect 16114 6780 16120 6792
rect 15694 6752 16120 6780
rect 15694 6749 15706 6752
rect 15648 6743 15706 6749
rect 1486 6672 1492 6724
rect 1544 6672 1550 6724
rect 15396 6712 15424 6743
rect 16114 6740 16120 6752
rect 16172 6780 16178 6792
rect 16942 6780 16948 6792
rect 16172 6752 16948 6780
rect 16172 6740 16178 6752
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 16574 6712 16580 6724
rect 15396 6684 16580 6712
rect 16574 6672 16580 6684
rect 16632 6672 16638 6724
rect 17052 6712 17080 6820
rect 17328 6780 17356 6820
rect 17880 6789 17908 6820
rect 17773 6783 17831 6789
rect 17773 6780 17785 6783
rect 17328 6752 17785 6780
rect 17773 6749 17785 6752
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6780 17923 6783
rect 18138 6780 18144 6792
rect 17911 6752 18144 6780
rect 17911 6749 17923 6752
rect 17865 6743 17923 6749
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 17221 6715 17279 6721
rect 17221 6712 17233 6715
rect 17052 6684 17233 6712
rect 17052 6656 17080 6684
rect 17221 6681 17233 6684
rect 17267 6681 17279 6715
rect 17221 6675 17279 6681
rect 17310 6672 17316 6724
rect 17368 6712 17374 6724
rect 17589 6715 17647 6721
rect 17589 6712 17601 6715
rect 17368 6684 17601 6712
rect 17368 6672 17374 6684
rect 17589 6681 17601 6684
rect 17635 6681 17647 6715
rect 17589 6675 17647 6681
rect 17954 6672 17960 6724
rect 18012 6672 18018 6724
rect 12894 6604 12900 6656
rect 12952 6604 12958 6656
rect 16761 6647 16819 6653
rect 16761 6613 16773 6647
rect 16807 6644 16819 6647
rect 17034 6644 17040 6656
rect 16807 6616 17040 6644
rect 16807 6613 16819 6616
rect 16761 6607 16819 6613
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17678 6644 17684 6656
rect 17175 6616 17684 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 17972 6644 18000 6672
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 17972 6616 18061 6644
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 18049 6607 18107 6613
rect 1104 6554 20792 6576
rect 1104 6502 7214 6554
rect 7266 6502 7278 6554
rect 7330 6502 7342 6554
rect 7394 6502 7406 6554
rect 7458 6502 7470 6554
rect 7522 6502 13214 6554
rect 13266 6502 13278 6554
rect 13330 6502 13342 6554
rect 13394 6502 13406 6554
rect 13458 6502 13470 6554
rect 13522 6502 19214 6554
rect 19266 6502 19278 6554
rect 19330 6502 19342 6554
rect 19394 6502 19406 6554
rect 19458 6502 19470 6554
rect 19522 6502 20792 6554
rect 1104 6480 20792 6502
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 7558 6440 7564 6452
rect 6328 6412 7564 6440
rect 6328 6400 6334 6412
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 9493 6443 9551 6449
rect 9493 6409 9505 6443
rect 9539 6440 9551 6443
rect 9582 6440 9588 6452
rect 9539 6412 9588 6440
rect 9539 6409 9551 6412
rect 9493 6403 9551 6409
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 12802 6440 12808 6452
rect 12360 6412 12808 6440
rect 6932 6344 8510 6372
rect 6932 6316 6960 6344
rect 2774 6264 2780 6316
rect 2832 6264 2838 6316
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2924 6276 3065 6304
rect 2924 6264 2930 6276
rect 3053 6273 3065 6276
rect 3099 6304 3111 6307
rect 3970 6304 3976 6316
rect 3099 6276 3976 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 6914 6264 6920 6316
rect 6972 6264 6978 6316
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 12360 6313 12388 6412
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 14093 6443 14151 6449
rect 12952 6412 13952 6440
rect 12952 6400 12958 6412
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7616 6276 7757 6304
rect 7616 6264 7622 6276
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 12345 6307 12403 6313
rect 12345 6304 12357 6307
rect 11011 6276 12357 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 12345 6273 12357 6276
rect 12391 6273 12403 6307
rect 12345 6267 12403 6273
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 13924 6304 13952 6412
rect 14093 6409 14105 6443
rect 14139 6409 14151 6443
rect 14093 6403 14151 6409
rect 14108 6372 14136 6403
rect 17034 6400 17040 6452
rect 17092 6400 17098 6452
rect 17678 6400 17684 6452
rect 17736 6440 17742 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 17736 6412 18061 6440
rect 17736 6400 17742 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 18138 6400 18144 6452
rect 18196 6400 18202 6452
rect 14461 6375 14519 6381
rect 14461 6372 14473 6375
rect 14108 6344 14473 6372
rect 14461 6341 14473 6344
rect 14507 6341 14519 6375
rect 14461 6335 14519 6341
rect 14185 6307 14243 6313
rect 14185 6304 14197 6307
rect 13924 6276 14197 6304
rect 14185 6273 14197 6276
rect 14231 6273 14243 6307
rect 16925 6307 16983 6313
rect 14185 6267 14243 6273
rect 8018 6196 8024 6248
rect 8076 6196 8082 6248
rect 11054 6196 11060 6248
rect 11112 6196 11118 6248
rect 12618 6196 12624 6248
rect 12676 6196 12682 6248
rect 13740 6236 13768 6264
rect 15580 6236 15608 6290
rect 16925 6273 16937 6307
rect 16971 6304 16983 6307
rect 17052 6304 17080 6400
rect 18156 6372 18184 6400
rect 18478 6375 18536 6381
rect 18478 6372 18490 6375
rect 18156 6344 18490 6372
rect 18478 6341 18490 6344
rect 18524 6341 18536 6375
rect 18478 6335 18536 6341
rect 16971 6276 17080 6304
rect 18233 6307 18291 6313
rect 16971 6273 16983 6276
rect 16925 6267 16983 6273
rect 18233 6273 18245 6307
rect 18279 6304 18291 6307
rect 18322 6304 18328 6316
rect 18279 6276 18328 6304
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 13740 6208 15608 6236
rect 16485 6239 16543 6245
rect 16485 6205 16497 6239
rect 16531 6236 16543 6239
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16531 6208 16681 6236
rect 16531 6205 16543 6208
rect 16485 6199 16543 6205
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 16669 6199 16727 6205
rect 2590 6060 2596 6112
rect 2648 6060 2654 6112
rect 3142 6060 3148 6112
rect 3200 6060 3206 6112
rect 10686 6060 10692 6112
rect 10744 6060 10750 6112
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 13044 6072 15945 6100
rect 13044 6060 13050 6072
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 15933 6063 15991 6069
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 16684 6100 16712 6199
rect 18138 6100 18144 6112
rect 16632 6072 18144 6100
rect 16632 6060 16638 6072
rect 18138 6060 18144 6072
rect 18196 6100 18202 6112
rect 18248 6100 18276 6267
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 18196 6072 18276 6100
rect 18196 6060 18202 6072
rect 19610 6060 19616 6112
rect 19668 6060 19674 6112
rect 1104 6010 20792 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 10214 6010
rect 10266 5958 10278 6010
rect 10330 5958 10342 6010
rect 10394 5958 10406 6010
rect 10458 5958 10470 6010
rect 10522 5958 16214 6010
rect 16266 5958 16278 6010
rect 16330 5958 16342 6010
rect 16394 5958 16406 6010
rect 16458 5958 16470 6010
rect 16522 5958 20792 6010
rect 1104 5936 20792 5958
rect 2130 5896 2136 5908
rect 1872 5868 2136 5896
rect 1872 5769 1900 5868
rect 2130 5856 2136 5868
rect 2188 5896 2194 5908
rect 2866 5896 2872 5908
rect 2188 5868 2872 5896
rect 2188 5856 2194 5868
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3142 5856 3148 5908
rect 3200 5856 3206 5908
rect 6089 5899 6147 5905
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6270 5896 6276 5908
rect 6135 5868 6276 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5729 1915 5763
rect 1857 5723 1915 5729
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5760 2191 5763
rect 2590 5760 2596 5772
rect 2179 5732 2596 5760
rect 2179 5729 2191 5732
rect 2133 5723 2191 5729
rect 2590 5720 2596 5732
rect 2648 5720 2654 5772
rect 3160 5760 3188 5856
rect 6196 5769 6224 5868
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 7929 5899 7987 5905
rect 7929 5865 7941 5899
rect 7975 5896 7987 5899
rect 8018 5896 8024 5908
rect 7975 5868 8024 5896
rect 7975 5865 7987 5868
rect 7929 5859 7987 5865
rect 8018 5856 8024 5868
rect 8076 5856 8082 5908
rect 11054 5856 11060 5908
rect 11112 5856 11118 5908
rect 12434 5856 12440 5908
rect 12492 5856 12498 5908
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 13081 5899 13139 5905
rect 13081 5896 13093 5899
rect 12676 5868 13093 5896
rect 12676 5856 12682 5868
rect 13081 5865 13093 5868
rect 13127 5865 13139 5899
rect 13081 5859 13139 5865
rect 16574 5856 16580 5908
rect 16632 5856 16638 5908
rect 16666 5856 16672 5908
rect 16724 5896 16730 5908
rect 16761 5899 16819 5905
rect 16761 5896 16773 5899
rect 16724 5868 16773 5896
rect 16724 5856 16730 5868
rect 16761 5865 16773 5868
rect 16807 5865 16819 5899
rect 16761 5859 16819 5865
rect 3605 5763 3663 5769
rect 3160 5732 3556 5760
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 3528 5692 3556 5732
rect 3605 5729 3617 5763
rect 3651 5760 3663 5763
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 3651 5732 4077 5760
rect 3651 5729 3663 5732
rect 3605 5723 3663 5729
rect 4065 5729 4077 5732
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 6181 5763 6239 5769
rect 6181 5729 6193 5763
rect 6227 5729 6239 5763
rect 6181 5723 6239 5729
rect 6822 5720 6828 5772
rect 6880 5760 6886 5772
rect 11072 5760 11100 5856
rect 11425 5831 11483 5837
rect 11425 5797 11437 5831
rect 11471 5828 11483 5831
rect 12802 5828 12808 5840
rect 11471 5800 12808 5828
rect 11471 5797 11483 5800
rect 11425 5791 11483 5797
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 11885 5763 11943 5769
rect 11885 5760 11897 5763
rect 6880 5732 8064 5760
rect 11072 5732 11897 5760
rect 6880 5720 6886 5732
rect 8036 5701 8064 5732
rect 11885 5729 11897 5732
rect 11931 5760 11943 5763
rect 12069 5763 12127 5769
rect 12069 5760 12081 5763
rect 11931 5732 12081 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 12069 5729 12081 5732
rect 12115 5729 12127 5763
rect 12069 5723 12127 5729
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3528 5664 3801 5692
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 8021 5695 8079 5701
rect 3789 5655 3847 5661
rect 3358 5596 4476 5624
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 2866 5556 2872 5568
rect 1627 5528 2872 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 4448 5556 4476 5596
rect 4798 5556 4804 5568
rect 4448 5528 4804 5556
rect 4798 5516 4804 5528
rect 4856 5556 4862 5568
rect 5074 5556 5080 5568
rect 4856 5528 5080 5556
rect 4856 5516 4862 5528
rect 5074 5516 5080 5528
rect 5132 5556 5138 5568
rect 5184 5556 5212 5678
rect 8021 5661 8033 5695
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5692 8723 5695
rect 9030 5692 9036 5704
rect 8711 5664 9036 5692
rect 8711 5661 8723 5664
rect 8665 5655 8723 5661
rect 5460 5596 6408 5624
rect 5460 5556 5488 5596
rect 5132 5528 5488 5556
rect 5132 5516 5138 5528
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 6380 5556 6408 5596
rect 6454 5584 6460 5636
rect 6512 5584 6518 5636
rect 6914 5624 6920 5636
rect 6656 5596 6920 5624
rect 6656 5556 6684 5596
rect 6914 5584 6920 5596
rect 6972 5584 6978 5636
rect 8496 5624 8524 5655
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 9508 5624 9536 5652
rect 8496 5596 9536 5624
rect 9784 5624 9812 5655
rect 10042 5652 10048 5704
rect 10100 5652 10106 5704
rect 10312 5695 10370 5701
rect 10312 5661 10324 5695
rect 10358 5692 10370 5695
rect 10686 5692 10692 5704
rect 10358 5664 10692 5692
rect 10358 5661 10370 5664
rect 10312 5655 10370 5661
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 11698 5652 11704 5704
rect 11756 5652 11762 5704
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 11517 5627 11575 5633
rect 11517 5624 11529 5627
rect 9784 5596 11529 5624
rect 11517 5593 11529 5596
rect 11563 5593 11575 5627
rect 11992 5624 12020 5655
rect 12158 5652 12164 5704
rect 12216 5652 12222 5704
rect 12618 5652 12624 5704
rect 12676 5652 12682 5704
rect 12820 5701 12848 5788
rect 18138 5720 18144 5772
rect 18196 5720 18202 5772
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 12986 5652 12992 5704
rect 13044 5652 13050 5704
rect 13078 5652 13084 5704
rect 13136 5692 13142 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 13136 5664 13277 5692
rect 13136 5652 13142 5664
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 13265 5655 13323 5661
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 11992 5596 12725 5624
rect 11517 5587 11575 5593
rect 12544 5568 12572 5596
rect 12713 5593 12725 5596
rect 12759 5593 12771 5627
rect 12713 5587 12771 5593
rect 17678 5584 17684 5636
rect 17736 5624 17742 5636
rect 17874 5627 17932 5633
rect 17874 5624 17886 5627
rect 17736 5596 17886 5624
rect 17736 5584 17742 5596
rect 17874 5593 17886 5596
rect 17920 5593 17932 5627
rect 17874 5587 17932 5593
rect 6380 5528 6684 5556
rect 8205 5559 8263 5565
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8478 5556 8484 5568
rect 8251 5528 8484 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 8570 5516 8576 5568
rect 8628 5516 8634 5568
rect 9950 5516 9956 5568
rect 10008 5516 10014 5568
rect 12526 5516 12532 5568
rect 12584 5516 12590 5568
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 13722 5556 13728 5568
rect 12676 5528 13728 5556
rect 12676 5516 12682 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 1104 5466 20792 5488
rect 1104 5414 7214 5466
rect 7266 5414 7278 5466
rect 7330 5414 7342 5466
rect 7394 5414 7406 5466
rect 7458 5414 7470 5466
rect 7522 5414 13214 5466
rect 13266 5414 13278 5466
rect 13330 5414 13342 5466
rect 13394 5414 13406 5466
rect 13458 5414 13470 5466
rect 13522 5414 19214 5466
rect 19266 5414 19278 5466
rect 19330 5414 19342 5466
rect 19394 5414 19406 5466
rect 19458 5414 19470 5466
rect 19522 5414 20792 5466
rect 1104 5392 20792 5414
rect 2774 5312 2780 5364
rect 2832 5312 2838 5364
rect 5534 5352 5540 5364
rect 3804 5324 5540 5352
rect 3237 5287 3295 5293
rect 3237 5253 3249 5287
rect 3283 5284 3295 5287
rect 3283 5256 3648 5284
rect 3283 5253 3295 5256
rect 3237 5247 3295 5253
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5185 3571 5219
rect 3513 5179 3571 5185
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 3528 5080 3556 5179
rect 3620 5148 3648 5256
rect 3804 5225 3832 5324
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 7926 5352 7932 5364
rect 6227 5324 6592 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 4065 5287 4123 5293
rect 4065 5284 4077 5287
rect 3896 5256 4077 5284
rect 3896 5228 3924 5256
rect 4065 5253 4077 5256
rect 4111 5253 4123 5287
rect 6270 5284 6276 5296
rect 5934 5256 6276 5284
rect 4065 5247 4123 5253
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 6564 5284 6592 5324
rect 7024 5324 7932 5352
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 6564 5256 6653 5284
rect 6641 5253 6653 5256
rect 6687 5253 6699 5287
rect 7024 5284 7052 5324
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 9326 5355 9384 5361
rect 9326 5321 9338 5355
rect 9372 5352 9384 5355
rect 10042 5352 10048 5364
rect 9372 5324 10048 5352
rect 9372 5321 9384 5324
rect 9326 5315 9384 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5321 11391 5355
rect 11333 5315 11391 5321
rect 11517 5355 11575 5361
rect 11517 5321 11529 5355
rect 11563 5352 11575 5355
rect 11698 5352 11704 5364
rect 11563 5324 11704 5352
rect 11563 5321 11575 5324
rect 11517 5315 11575 5321
rect 7098 5284 7104 5296
rect 7024 5256 7104 5284
rect 6641 5247 6699 5253
rect 7098 5244 7104 5256
rect 7156 5244 7162 5296
rect 8478 5244 8484 5296
rect 8536 5284 8542 5296
rect 8536 5256 9220 5284
rect 8536 5244 8542 5256
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5216 3755 5219
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3743 5188 3801 5216
rect 3743 5185 3755 5188
rect 3697 5179 3755 5185
rect 3789 5185 3801 5188
rect 3835 5185 3847 5219
rect 3789 5179 3847 5185
rect 3878 5176 3884 5228
rect 3936 5176 3942 5228
rect 3970 5176 3976 5228
rect 4028 5176 4034 5228
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4172 5148 4200 5179
rect 8570 5176 8576 5228
rect 8628 5176 8634 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8680 5188 8769 5216
rect 4433 5151 4491 5157
rect 4433 5148 4445 5151
rect 3620 5120 4200 5148
rect 2924 5052 3556 5080
rect 2924 5040 2930 5052
rect 3510 4972 3516 5024
rect 3568 4972 3574 5024
rect 4172 5012 4200 5120
rect 4356 5120 4445 5148
rect 4356 5089 4384 5120
rect 4433 5117 4445 5120
rect 4479 5117 4491 5151
rect 4433 5111 4491 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4755 5120 6316 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4341 5083 4399 5089
rect 4341 5049 4353 5083
rect 4387 5049 4399 5083
rect 6288 5080 6316 5120
rect 6362 5108 6368 5160
rect 6420 5108 6426 5160
rect 8588 5148 8616 5176
rect 6472 5120 8616 5148
rect 6472 5080 6500 5120
rect 6288 5052 6500 5080
rect 8113 5083 8171 5089
rect 4341 5043 4399 5049
rect 8113 5049 8125 5083
rect 8159 5080 8171 5083
rect 8202 5080 8208 5092
rect 8159 5052 8208 5080
rect 8159 5049 8171 5052
rect 8113 5043 8171 5049
rect 8202 5040 8208 5052
rect 8260 5080 8266 5092
rect 8680 5080 8708 5188
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 8260 5052 8708 5080
rect 8260 5040 8266 5052
rect 4798 5012 4804 5024
rect 4172 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 8956 5012 8984 5179
rect 9030 5176 9036 5228
rect 9088 5176 9094 5228
rect 9192 5225 9220 5256
rect 9490 5244 9496 5296
rect 9548 5284 9554 5296
rect 9585 5287 9643 5293
rect 9585 5284 9597 5287
rect 9548 5256 9597 5284
rect 9548 5244 9554 5256
rect 9585 5253 9597 5256
rect 9631 5253 9643 5287
rect 9585 5247 9643 5253
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 10198 5287 10256 5293
rect 10198 5284 10210 5287
rect 10008 5256 10210 5284
rect 10008 5244 10014 5256
rect 10198 5253 10210 5256
rect 10244 5253 10256 5287
rect 11348 5284 11376 5315
rect 11698 5312 11704 5324
rect 11756 5312 11762 5364
rect 12805 5355 12863 5361
rect 12805 5321 12817 5355
rect 12851 5352 12863 5355
rect 13078 5352 13084 5364
rect 12851 5324 13084 5352
rect 12851 5321 12863 5324
rect 12805 5315 12863 5321
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 18049 5355 18107 5361
rect 14568 5324 15148 5352
rect 12526 5284 12532 5296
rect 11348 5256 12532 5284
rect 10198 5247 10256 5253
rect 9171 5219 9229 5225
rect 9171 5185 9183 5219
rect 9217 5216 9229 5219
rect 9398 5216 9404 5228
rect 9217 5188 9404 5216
rect 9217 5185 9229 5188
rect 9171 5179 9229 5185
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 9674 5176 9680 5228
rect 9732 5176 9738 5228
rect 11716 5225 11744 5256
rect 12526 5244 12532 5256
rect 12584 5284 12590 5296
rect 14458 5284 14464 5296
rect 12584 5256 12940 5284
rect 14398 5256 14464 5284
rect 12584 5244 12590 5256
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 12158 5216 12164 5228
rect 11931 5188 12164 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12618 5176 12624 5228
rect 12676 5176 12682 5228
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9508 5120 9965 5148
rect 9508 5024 9536 5120
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 12636 5148 12664 5176
rect 12912 5157 12940 5256
rect 14458 5244 14464 5256
rect 14516 5284 14522 5296
rect 14568 5284 14596 5324
rect 14516 5256 14596 5284
rect 15120 5284 15148 5324
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 18138 5352 18144 5364
rect 18095 5324 18144 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 18233 5355 18291 5361
rect 18233 5321 18245 5355
rect 18279 5352 18291 5355
rect 19702 5352 19708 5364
rect 18279 5324 19708 5352
rect 18279 5321 18291 5324
rect 18233 5315 18291 5321
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 15120 5256 15502 5284
rect 14516 5244 14522 5256
rect 18156 5216 18184 5312
rect 19368 5287 19426 5293
rect 19368 5253 19380 5287
rect 19414 5284 19426 5287
rect 19610 5284 19616 5296
rect 19414 5256 19616 5284
rect 19414 5253 19426 5256
rect 19368 5247 19426 5253
rect 19610 5244 19616 5256
rect 19668 5244 19674 5296
rect 20441 5219 20499 5225
rect 18156 5188 19656 5216
rect 12391 5120 12664 5148
rect 12897 5151 12955 5157
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 12897 5117 12909 5151
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 12618 5040 12624 5092
rect 12676 5040 12682 5092
rect 9122 5012 9128 5024
rect 6512 4984 9128 5012
rect 6512 4972 6518 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9490 4972 9496 5024
rect 9548 4972 9554 5024
rect 12912 5012 12940 5111
rect 13170 5108 13176 5160
rect 13228 5108 13234 5160
rect 14734 5108 14740 5160
rect 14792 5108 14798 5160
rect 19628 5157 19656 5188
rect 20441 5185 20453 5219
rect 20487 5216 20499 5219
rect 20806 5216 20812 5228
rect 20487 5188 20812 5216
rect 20487 5185 20499 5188
rect 20441 5179 20499 5185
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14844 5120 15025 5148
rect 14645 5083 14703 5089
rect 14645 5049 14657 5083
rect 14691 5080 14703 5083
rect 14844 5080 14872 5120
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15013 5111 15071 5117
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5117 19671 5151
rect 19613 5111 19671 5117
rect 14691 5052 14872 5080
rect 14691 5049 14703 5052
rect 14645 5043 14703 5049
rect 13354 5012 13360 5024
rect 12912 4984 13360 5012
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13722 4972 13728 5024
rect 13780 5012 13786 5024
rect 16485 5015 16543 5021
rect 16485 5012 16497 5015
rect 13780 4984 16497 5012
rect 13780 4972 13786 4984
rect 16485 4981 16497 4984
rect 16531 4981 16543 5015
rect 16485 4975 16543 4981
rect 20254 4972 20260 5024
rect 20312 4972 20318 5024
rect 1104 4922 20792 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 10214 4922
rect 10266 4870 10278 4922
rect 10330 4870 10342 4922
rect 10394 4870 10406 4922
rect 10458 4870 10470 4922
rect 10522 4870 16214 4922
rect 16266 4870 16278 4922
rect 16330 4870 16342 4922
rect 16394 4870 16406 4922
rect 16458 4870 16470 4922
rect 16522 4870 20792 4922
rect 1104 4848 20792 4870
rect 5534 4768 5540 4820
rect 5592 4768 5598 4820
rect 6273 4811 6331 4817
rect 6273 4777 6285 4811
rect 6319 4808 6331 4811
rect 6362 4808 6368 4820
rect 6319 4780 6368 4808
rect 6319 4777 6331 4780
rect 6273 4771 6331 4777
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 9490 4768 9496 4820
rect 9548 4768 9554 4820
rect 13081 4811 13139 4817
rect 13081 4777 13093 4811
rect 13127 4808 13139 4811
rect 13170 4808 13176 4820
rect 13127 4780 13176 4808
rect 13127 4777 13139 4780
rect 13081 4771 13139 4777
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13449 4811 13507 4817
rect 13449 4777 13461 4811
rect 13495 4808 13507 4811
rect 14734 4808 14740 4820
rect 13495 4780 14740 4808
rect 13495 4777 13507 4780
rect 13449 4771 13507 4777
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 5552 4672 5580 4768
rect 14369 4743 14427 4749
rect 14369 4709 14381 4743
rect 14415 4740 14427 4743
rect 14458 4740 14464 4752
rect 14415 4712 14464 4740
rect 14415 4709 14427 4712
rect 14369 4703 14427 4709
rect 14458 4700 14464 4712
rect 14516 4700 14522 4752
rect 4448 4644 5580 4672
rect 5721 4675 5779 4681
rect 4448 4613 4476 4644
rect 5721 4641 5733 4675
rect 5767 4672 5779 4675
rect 6454 4672 6460 4684
rect 5767 4644 6460 4672
rect 5767 4641 5779 4644
rect 5721 4635 5779 4641
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 5994 4604 6000 4616
rect 4856 4576 6000 4604
rect 4856 4564 4862 4576
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6196 4613 6224 4644
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8260 4576 8953 4604
rect 8260 4564 8266 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9214 4604 9220 4616
rect 9088 4576 9220 4604
rect 9088 4564 9094 4576
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9398 4613 9404 4616
rect 9355 4607 9404 4613
rect 9355 4573 9367 4607
rect 9401 4573 9404 4607
rect 9355 4567 9404 4573
rect 9398 4564 9404 4567
rect 9456 4564 9462 4616
rect 12897 4607 12955 4613
rect 12897 4573 12909 4607
rect 12943 4604 12955 4607
rect 12986 4604 12992 4616
rect 12943 4576 12992 4604
rect 12943 4573 12955 4576
rect 12897 4567 12955 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13078 4564 13084 4616
rect 13136 4564 13142 4616
rect 13354 4564 13360 4616
rect 13412 4564 13418 4616
rect 20254 4604 20260 4616
rect 14108 4576 20260 4604
rect 3878 4496 3884 4548
rect 3936 4496 3942 4548
rect 3970 4496 3976 4548
rect 4028 4536 4034 4548
rect 4617 4539 4675 4545
rect 4617 4536 4629 4539
rect 4028 4508 4629 4536
rect 4028 4496 4034 4508
rect 4617 4505 4629 4508
rect 4663 4505 4675 4539
rect 4617 4499 4675 4505
rect 4709 4539 4767 4545
rect 4709 4505 4721 4539
rect 4755 4505 4767 4539
rect 4709 4499 4767 4505
rect 5537 4539 5595 4545
rect 5537 4505 5549 4539
rect 5583 4505 5595 4539
rect 5537 4499 5595 4505
rect 3896 4468 3924 4496
rect 4724 4468 4752 4499
rect 3896 4440 4752 4468
rect 4985 4471 5043 4477
rect 4985 4437 4997 4471
rect 5031 4468 5043 4471
rect 5552 4468 5580 4499
rect 9122 4496 9128 4548
rect 9180 4496 9186 4548
rect 9674 4496 9680 4548
rect 9732 4536 9738 4548
rect 14108 4536 14136 4576
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 9732 4508 14136 4536
rect 9732 4496 9738 4508
rect 14182 4496 14188 4548
rect 14240 4496 14246 4548
rect 5031 4440 5580 4468
rect 9140 4468 9168 4496
rect 9950 4468 9956 4480
rect 9140 4440 9956 4468
rect 5031 4437 5043 4440
rect 4985 4431 5043 4437
rect 9950 4428 9956 4440
rect 10008 4428 10014 4480
rect 1104 4378 20792 4400
rect 1104 4326 7214 4378
rect 7266 4326 7278 4378
rect 7330 4326 7342 4378
rect 7394 4326 7406 4378
rect 7458 4326 7470 4378
rect 7522 4326 13214 4378
rect 13266 4326 13278 4378
rect 13330 4326 13342 4378
rect 13394 4326 13406 4378
rect 13458 4326 13470 4378
rect 13522 4326 19214 4378
rect 19266 4326 19278 4378
rect 19330 4326 19342 4378
rect 19394 4326 19406 4378
rect 19458 4326 19470 4378
rect 19522 4326 20792 4378
rect 1104 4304 20792 4326
rect 8202 4224 8208 4276
rect 8260 4264 8266 4276
rect 8260 4236 9536 4264
rect 8260 4224 8266 4236
rect 8220 4196 8248 4224
rect 7852 4168 8248 4196
rect 14 4088 20 4140
rect 72 4128 78 4140
rect 1486 4128 1492 4140
rect 72 4100 1492 4128
rect 72 4088 78 4100
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 7650 4088 7656 4140
rect 7708 4088 7714 4140
rect 7852 4137 7880 4168
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 9508 4128 9536 4236
rect 12158 4224 12164 4276
rect 12216 4224 12222 4276
rect 9876 4168 10180 4196
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9508 4100 9781 4128
rect 9769 4097 9781 4100
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 7926 4020 7932 4072
rect 7984 4020 7990 4072
rect 8202 4020 8208 4072
rect 8260 4020 8266 4072
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9398 4060 9404 4072
rect 8720 4032 9404 4060
rect 8720 4020 8726 4032
rect 9398 4020 9404 4032
rect 9456 4060 9462 4072
rect 9876 4060 9904 4168
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10152 4137 10180 4168
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10142 4131 10200 4137
rect 10142 4097 10154 4131
rect 10188 4097 10200 4131
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10142 4091 10200 4097
rect 10244 4100 10701 4128
rect 9456 4032 9904 4060
rect 9456 4020 9462 4032
rect 10060 3992 10088 4091
rect 9692 3964 10088 3992
rect 7650 3884 7656 3936
rect 7708 3884 7714 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9692 3933 9720 3964
rect 9677 3927 9735 3933
rect 9677 3924 9689 3927
rect 9272 3896 9689 3924
rect 9272 3884 9278 3896
rect 9677 3893 9689 3896
rect 9723 3893 9735 3927
rect 9677 3887 9735 3893
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 10244 3924 10272 4100
rect 10689 4097 10701 4100
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 12176 4128 12204 4224
rect 12618 4196 12624 4208
rect 12406 4168 12624 4196
rect 12406 4128 12434 4168
rect 12618 4156 12624 4168
rect 12676 4196 12682 4208
rect 12676 4168 12848 4196
rect 12676 4156 12682 4168
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 11747 4100 12204 4128
rect 12360 4100 12541 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 11974 4020 11980 4072
rect 12032 4020 12038 4072
rect 10321 3995 10379 4001
rect 10321 3961 10333 3995
rect 10367 3992 10379 3995
rect 10686 3992 10692 4004
rect 10367 3964 10692 3992
rect 10367 3961 10379 3964
rect 10321 3955 10379 3961
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 12360 4001 12388 4100
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4097 12771 4131
rect 12820 4128 12848 4168
rect 13078 4128 13084 4140
rect 12820 4100 13084 4128
rect 12713 4091 12771 4097
rect 12345 3995 12403 4001
rect 12345 3961 12357 3995
rect 12391 3961 12403 3995
rect 12345 3955 12403 3961
rect 12728 3936 12756 4091
rect 13078 4088 13084 4100
rect 13136 4128 13142 4140
rect 13136 4100 20668 4128
rect 13136 4088 13142 4100
rect 20640 4072 20668 4100
rect 20622 4020 20628 4072
rect 20680 4020 20686 4072
rect 10008 3896 10272 3924
rect 10008 3884 10014 3896
rect 10594 3884 10600 3936
rect 10652 3884 10658 3936
rect 11609 3927 11667 3933
rect 11609 3893 11621 3927
rect 11655 3924 11667 3927
rect 11882 3924 11888 3936
rect 11655 3896 11888 3924
rect 11655 3893 11667 3896
rect 11609 3887 11667 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12434 3884 12440 3936
rect 12492 3884 12498 3936
rect 12526 3884 12532 3936
rect 12584 3884 12590 3936
rect 12710 3884 12716 3936
rect 12768 3884 12774 3936
rect 1104 3834 20792 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 10214 3834
rect 10266 3782 10278 3834
rect 10330 3782 10342 3834
rect 10394 3782 10406 3834
rect 10458 3782 10470 3834
rect 10522 3782 16214 3834
rect 16266 3782 16278 3834
rect 16330 3782 16342 3834
rect 16394 3782 16406 3834
rect 16458 3782 16470 3834
rect 16522 3782 20792 3834
rect 1104 3760 20792 3782
rect 5994 3680 6000 3732
rect 6052 3680 6058 3732
rect 7180 3723 7238 3729
rect 7180 3689 7192 3723
rect 7226 3720 7238 3723
rect 7650 3720 7656 3732
rect 7226 3692 7656 3720
rect 7226 3689 7238 3692
rect 7180 3683 7238 3689
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 8202 3680 8208 3732
rect 8260 3720 8266 3732
rect 8665 3723 8723 3729
rect 8665 3720 8677 3723
rect 8260 3692 8677 3720
rect 8260 3680 8266 3692
rect 8665 3689 8677 3692
rect 8711 3689 8723 3723
rect 8665 3683 8723 3689
rect 9950 3680 9956 3732
rect 10008 3680 10014 3732
rect 10594 3720 10600 3732
rect 10244 3692 10600 3720
rect 9493 3655 9551 3661
rect 9493 3621 9505 3655
rect 9539 3621 9551 3655
rect 9493 3615 9551 3621
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3896 3488 3985 3516
rect 3896 3460 3924 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3516 4123 3519
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 4111 3488 4261 3516
rect 4111 3485 4123 3488
rect 4065 3479 4123 3485
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 6914 3476 6920 3528
rect 6972 3476 6978 3528
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 9398 3525 9404 3528
rect 8941 3519 8999 3525
rect 8941 3485 8953 3519
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 9355 3519 9404 3525
rect 9355 3485 9367 3519
rect 9401 3485 9404 3519
rect 9355 3479 9404 3485
rect 3878 3408 3884 3460
rect 3936 3408 3942 3460
rect 4522 3408 4528 3460
rect 4580 3408 4586 3460
rect 5074 3408 5080 3460
rect 5132 3408 5138 3460
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8956 3380 8984 3479
rect 9398 3476 9404 3479
rect 9456 3476 9462 3528
rect 9508 3516 9536 3615
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3584 10195 3587
rect 10244 3584 10272 3692
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 11882 3680 11888 3732
rect 11940 3680 11946 3732
rect 10183 3556 10272 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10410 3544 10416 3596
rect 10468 3544 10474 3596
rect 11900 3584 11928 3680
rect 11900 3556 12112 3584
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9508 3488 9781 3516
rect 9769 3485 9781 3488
rect 9815 3485 9827 3519
rect 11974 3516 11980 3528
rect 9769 3479 9827 3485
rect 11716 3488 11980 3516
rect 9122 3408 9128 3460
rect 9180 3408 9186 3460
rect 9214 3408 9220 3460
rect 9272 3408 9278 3460
rect 9324 3420 10902 3448
rect 9324 3392 9352 3420
rect 8168 3352 8984 3380
rect 8168 3340 8174 3352
rect 9306 3340 9312 3392
rect 9364 3340 9370 3392
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 11716 3380 11744 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12084 3516 12112 3556
rect 12233 3519 12291 3525
rect 12233 3516 12245 3519
rect 12084 3488 12245 3516
rect 12233 3485 12245 3488
rect 12279 3485 12291 3519
rect 12526 3516 12532 3528
rect 12233 3479 12291 3485
rect 12406 3488 12532 3516
rect 12406 3448 12434 3488
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 11808 3420 12434 3448
rect 11808 3392 11836 3420
rect 10008 3352 11744 3380
rect 10008 3340 10014 3352
rect 11790 3340 11796 3392
rect 11848 3340 11854 3392
rect 11882 3340 11888 3392
rect 11940 3340 11946 3392
rect 12342 3340 12348 3392
rect 12400 3380 12406 3392
rect 12526 3380 12532 3392
rect 12400 3352 12532 3380
rect 12400 3340 12406 3352
rect 12526 3340 12532 3352
rect 12584 3380 12590 3392
rect 13357 3383 13415 3389
rect 13357 3380 13369 3383
rect 12584 3352 13369 3380
rect 12584 3340 12590 3352
rect 13357 3349 13369 3352
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 1104 3290 20792 3312
rect 1104 3238 7214 3290
rect 7266 3238 7278 3290
rect 7330 3238 7342 3290
rect 7394 3238 7406 3290
rect 7458 3238 7470 3290
rect 7522 3238 13214 3290
rect 13266 3238 13278 3290
rect 13330 3238 13342 3290
rect 13394 3238 13406 3290
rect 13458 3238 13470 3290
rect 13522 3238 19214 3290
rect 19266 3238 19278 3290
rect 19330 3238 19342 3290
rect 19394 3238 19406 3290
rect 19458 3238 19470 3290
rect 19522 3238 20792 3290
rect 1104 3216 20792 3238
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 4580 3148 5273 3176
rect 4580 3136 4586 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5261 3139 5319 3145
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 7926 3176 7932 3188
rect 7883 3148 7932 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 8941 3179 8999 3185
rect 8941 3145 8953 3179
rect 8987 3176 8999 3179
rect 10410 3176 10416 3188
rect 8987 3148 10416 3176
rect 8987 3145 8999 3148
rect 8941 3139 8999 3145
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 10686 3136 10692 3188
rect 10744 3136 10750 3188
rect 11790 3176 11796 3188
rect 11624 3148 11796 3176
rect 3510 3068 3516 3120
rect 3568 3108 3574 3120
rect 3789 3111 3847 3117
rect 3789 3108 3801 3111
rect 3568 3080 3801 3108
rect 3568 3068 3574 3080
rect 3789 3077 3801 3080
rect 3835 3077 3847 3111
rect 5074 3108 5080 3120
rect 5014 3080 5080 3108
rect 3789 3071 3847 3077
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 6932 3040 6960 3136
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 6932 3012 7757 3040
rect 7745 3009 7757 3012
rect 7791 3040 7803 3043
rect 8662 3040 8668 3052
rect 7791 3012 8668 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9306 3000 9312 3052
rect 9364 3000 9370 3052
rect 10704 3049 10732 3136
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 3878 2972 3884 2984
rect 3559 2944 3884 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 3878 2932 3884 2944
rect 3936 2972 3942 2984
rect 9674 2972 9680 2984
rect 3936 2944 9680 2972
rect 3936 2932 3942 2944
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 10413 2975 10471 2981
rect 10413 2941 10425 2975
rect 10459 2972 10471 2975
rect 11624 2972 11652 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11974 3136 11980 3188
rect 12032 3136 12038 3188
rect 12066 3136 12072 3188
rect 12124 3136 12130 3188
rect 14550 3176 14556 3188
rect 14016 3148 14556 3176
rect 11790 3049 11796 3052
rect 11788 3040 11796 3049
rect 11751 3012 11796 3040
rect 11788 3003 11796 3012
rect 11790 3000 11796 3003
rect 11848 3000 11854 3052
rect 11992 3049 12020 3136
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3009 12035 3043
rect 12084 3040 12112 3136
rect 12526 3108 12532 3120
rect 12360 3080 12532 3108
rect 12360 3049 12388 3080
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 14016 3108 14044 3148
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 13846 3080 14044 3108
rect 14568 3108 14596 3136
rect 14918 3108 14924 3120
rect 14568 3080 14924 3108
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 12161 3043 12219 3049
rect 12161 3040 12173 3043
rect 12084 3012 12173 3040
rect 11977 3003 12035 3009
rect 12161 3009 12173 3012
rect 12207 3009 12219 3043
rect 12161 3003 12219 3009
rect 12345 3043 12403 3049
rect 12345 3009 12357 3043
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 10459 2944 11652 2972
rect 10459 2941 10471 2944
rect 10413 2935 10471 2941
rect 11606 2864 11612 2916
rect 11664 2864 11670 2916
rect 11900 2836 11928 3003
rect 12618 2932 12624 2984
rect 12676 2932 12682 2984
rect 14182 2932 14188 2984
rect 14240 2932 14246 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 14292 2944 14473 2972
rect 14093 2907 14151 2913
rect 14093 2873 14105 2907
rect 14139 2904 14151 2907
rect 14292 2904 14320 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 14139 2876 14320 2904
rect 14139 2873 14151 2876
rect 14093 2867 14151 2873
rect 12710 2836 12716 2848
rect 11900 2808 12716 2836
rect 12710 2796 12716 2808
rect 12768 2836 12774 2848
rect 15933 2839 15991 2845
rect 15933 2836 15945 2839
rect 12768 2808 15945 2836
rect 12768 2796 12774 2808
rect 15933 2805 15945 2808
rect 15979 2805 15991 2839
rect 15933 2799 15991 2805
rect 1104 2746 20792 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 10214 2746
rect 10266 2694 10278 2746
rect 10330 2694 10342 2746
rect 10394 2694 10406 2746
rect 10458 2694 10470 2746
rect 10522 2694 16214 2746
rect 16266 2694 16278 2746
rect 16330 2694 16342 2746
rect 16394 2694 16406 2746
rect 16458 2694 16470 2746
rect 16522 2694 20792 2746
rect 1104 2672 20792 2694
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 8754 2632 8760 2644
rect 5491 2604 8760 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 12618 2592 12624 2644
rect 12676 2592 12682 2644
rect 12897 2635 12955 2641
rect 12897 2601 12909 2635
rect 12943 2632 12955 2635
rect 14182 2632 14188 2644
rect 12943 2604 14188 2632
rect 12943 2601 12955 2604
rect 12897 2595 12955 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 9732 2468 10701 2496
rect 9732 2456 9738 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 10410 2388 10416 2440
rect 10468 2388 10474 2440
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12584 2400 12817 2428
rect 12584 2388 12590 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 15194 2388 15200 2440
rect 15252 2428 15258 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15252 2400 15761 2428
rect 15252 2388 15258 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 15562 2320 15568 2372
rect 15620 2320 15626 2372
rect 1104 2202 20792 2224
rect 1104 2150 7214 2202
rect 7266 2150 7278 2202
rect 7330 2150 7342 2202
rect 7394 2150 7406 2202
rect 7458 2150 7470 2202
rect 7522 2150 13214 2202
rect 13266 2150 13278 2202
rect 13330 2150 13342 2202
rect 13394 2150 13406 2202
rect 13458 2150 13470 2202
rect 13522 2150 19214 2202
rect 19266 2150 19278 2202
rect 19330 2150 19342 2202
rect 19394 2150 19406 2202
rect 19458 2150 19470 2202
rect 19522 2150 20792 2202
rect 1104 2128 20792 2150
<< via1 >>
rect 7214 21734 7266 21786
rect 7278 21734 7330 21786
rect 7342 21734 7394 21786
rect 7406 21734 7458 21786
rect 7470 21734 7522 21786
rect 13214 21734 13266 21786
rect 13278 21734 13330 21786
rect 13342 21734 13394 21786
rect 13406 21734 13458 21786
rect 13470 21734 13522 21786
rect 19214 21734 19266 21786
rect 19278 21734 19330 21786
rect 19342 21734 19394 21786
rect 19406 21734 19458 21786
rect 19470 21734 19522 21786
rect 3332 21539 3384 21548
rect 3332 21505 3341 21539
rect 3341 21505 3375 21539
rect 3375 21505 3384 21539
rect 3332 21496 3384 21505
rect 13820 21496 13872 21548
rect 17776 21539 17828 21548
rect 17776 21505 17785 21539
rect 17785 21505 17819 21539
rect 17819 21505 17828 21539
rect 17776 21496 17828 21505
rect 18144 21496 18196 21548
rect 18696 21496 18748 21548
rect 20260 21539 20312 21548
rect 20260 21505 20269 21539
rect 20269 21505 20303 21539
rect 20303 21505 20312 21539
rect 20260 21496 20312 21505
rect 14372 21471 14424 21480
rect 14372 21437 14381 21471
rect 14381 21437 14415 21471
rect 14415 21437 14424 21471
rect 14372 21428 14424 21437
rect 17960 21471 18012 21480
rect 17960 21437 17969 21471
rect 17969 21437 18003 21471
rect 18003 21437 18012 21471
rect 17960 21428 18012 21437
rect 4804 21292 4856 21344
rect 12440 21292 12492 21344
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 18236 21335 18288 21344
rect 18236 21301 18245 21335
rect 18245 21301 18279 21335
rect 18279 21301 18288 21335
rect 18236 21292 18288 21301
rect 18328 21292 18380 21344
rect 18604 21292 18656 21344
rect 20444 21292 20496 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 10214 21190 10266 21242
rect 10278 21190 10330 21242
rect 10342 21190 10394 21242
rect 10406 21190 10458 21242
rect 10470 21190 10522 21242
rect 16214 21190 16266 21242
rect 16278 21190 16330 21242
rect 16342 21190 16394 21242
rect 16406 21190 16458 21242
rect 16470 21190 16522 21242
rect 7012 20884 7064 20936
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 8392 20884 8444 20936
rect 4896 20791 4948 20800
rect 4896 20757 4905 20791
rect 4905 20757 4939 20791
rect 4939 20757 4948 20791
rect 4896 20748 4948 20757
rect 7564 20791 7616 20800
rect 7564 20757 7573 20791
rect 7573 20757 7607 20791
rect 7607 20757 7616 20791
rect 7564 20748 7616 20757
rect 8300 20748 8352 20800
rect 12440 21088 12492 21140
rect 14372 21088 14424 21140
rect 18052 21088 18104 21140
rect 18788 21088 18840 21140
rect 12624 20884 12676 20936
rect 8760 20816 8812 20868
rect 11612 20816 11664 20868
rect 15476 20884 15528 20936
rect 15568 20927 15620 20936
rect 15568 20893 15577 20927
rect 15577 20893 15611 20927
rect 15611 20893 15620 20927
rect 15568 20884 15620 20893
rect 17316 20927 17368 20936
rect 17316 20893 17325 20927
rect 17325 20893 17359 20927
rect 17359 20893 17368 20927
rect 17316 20884 17368 20893
rect 15200 20816 15252 20868
rect 17960 20816 18012 20868
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 10324 20748 10376 20757
rect 10784 20791 10836 20800
rect 10784 20757 10793 20791
rect 10793 20757 10827 20791
rect 10827 20757 10836 20791
rect 10784 20748 10836 20757
rect 12532 20791 12584 20800
rect 12532 20757 12541 20791
rect 12541 20757 12575 20791
rect 12575 20757 12584 20791
rect 12532 20748 12584 20757
rect 14188 20791 14240 20800
rect 14188 20757 14197 20791
rect 14197 20757 14231 20791
rect 14231 20757 14240 20791
rect 14188 20748 14240 20757
rect 7214 20646 7266 20698
rect 7278 20646 7330 20698
rect 7342 20646 7394 20698
rect 7406 20646 7458 20698
rect 7470 20646 7522 20698
rect 13214 20646 13266 20698
rect 13278 20646 13330 20698
rect 13342 20646 13394 20698
rect 13406 20646 13458 20698
rect 13470 20646 13522 20698
rect 19214 20646 19266 20698
rect 19278 20646 19330 20698
rect 19342 20646 19394 20698
rect 19406 20646 19458 20698
rect 19470 20646 19522 20698
rect 8760 20544 8812 20596
rect 11612 20587 11664 20596
rect 11612 20553 11621 20587
rect 11621 20553 11655 20587
rect 11655 20553 11664 20587
rect 11612 20544 11664 20553
rect 7564 20519 7616 20528
rect 7564 20485 7582 20519
rect 7582 20485 7616 20519
rect 7564 20476 7616 20485
rect 10876 20476 10928 20528
rect 12440 20476 12492 20528
rect 12532 20476 12584 20528
rect 14188 20476 14240 20528
rect 4896 20451 4948 20460
rect 4896 20417 4905 20451
rect 4905 20417 4939 20451
rect 4939 20417 4948 20451
rect 4896 20408 4948 20417
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 4068 20204 4120 20256
rect 5816 20247 5868 20256
rect 5816 20213 5825 20247
rect 5825 20213 5859 20247
rect 5859 20213 5868 20247
rect 5816 20204 5868 20213
rect 7012 20408 7064 20460
rect 10140 20408 10192 20460
rect 10324 20408 10376 20460
rect 8300 20340 8352 20392
rect 6552 20204 6604 20256
rect 13728 20408 13780 20460
rect 16948 20519 17000 20528
rect 16948 20485 16982 20519
rect 16982 20485 17000 20519
rect 16948 20476 17000 20485
rect 17776 20476 17828 20528
rect 18144 20476 18196 20528
rect 17316 20408 17368 20460
rect 18328 20408 18380 20460
rect 12624 20204 12676 20256
rect 15016 20247 15068 20256
rect 15016 20213 15025 20247
rect 15025 20213 15059 20247
rect 15059 20213 15068 20247
rect 15016 20204 15068 20213
rect 15200 20204 15252 20256
rect 15568 20204 15620 20256
rect 17960 20204 18012 20256
rect 19616 20247 19668 20256
rect 19616 20213 19625 20247
rect 19625 20213 19659 20247
rect 19659 20213 19668 20247
rect 19616 20204 19668 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 10214 20102 10266 20154
rect 10278 20102 10330 20154
rect 10342 20102 10394 20154
rect 10406 20102 10458 20154
rect 10470 20102 10522 20154
rect 16214 20102 16266 20154
rect 16278 20102 16330 20154
rect 16342 20102 16394 20154
rect 16406 20102 16458 20154
rect 16470 20102 16522 20154
rect 7104 20000 7156 20052
rect 10140 20000 10192 20052
rect 12624 20000 12676 20052
rect 12900 20043 12952 20052
rect 12900 20009 12909 20043
rect 12909 20009 12943 20043
rect 12943 20009 12952 20043
rect 12900 20000 12952 20009
rect 15200 20000 15252 20052
rect 16948 20043 17000 20052
rect 16948 20009 16957 20043
rect 16957 20009 16991 20043
rect 16991 20009 17000 20043
rect 16948 20000 17000 20009
rect 17316 20000 17368 20052
rect 18144 20000 18196 20052
rect 18328 20000 18380 20052
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 6000 19796 6052 19848
rect 6276 19839 6328 19848
rect 6276 19805 6285 19839
rect 6285 19805 6319 19839
rect 6319 19805 6328 19839
rect 6276 19796 6328 19805
rect 6460 19839 6512 19848
rect 6460 19805 6469 19839
rect 6469 19805 6503 19839
rect 6503 19805 6512 19839
rect 6460 19796 6512 19805
rect 6552 19796 6604 19848
rect 10784 19839 10836 19848
rect 10784 19805 10818 19839
rect 10818 19805 10836 19839
rect 10784 19796 10836 19805
rect 11796 19728 11848 19780
rect 12440 19796 12492 19848
rect 13728 19796 13780 19848
rect 4068 19703 4120 19712
rect 4068 19669 4077 19703
rect 4077 19669 4111 19703
rect 4111 19669 4120 19703
rect 4068 19660 4120 19669
rect 6368 19703 6420 19712
rect 6368 19669 6377 19703
rect 6377 19669 6411 19703
rect 6411 19669 6420 19703
rect 6368 19660 6420 19669
rect 11152 19660 11204 19712
rect 12256 19703 12308 19712
rect 12256 19669 12265 19703
rect 12265 19669 12299 19703
rect 12299 19669 12308 19703
rect 12256 19660 12308 19669
rect 13820 19728 13872 19780
rect 14188 19796 14240 19848
rect 15568 19839 15620 19848
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 18788 19839 18840 19848
rect 18788 19805 18806 19839
rect 18806 19805 18840 19839
rect 18788 19796 18840 19805
rect 16120 19728 16172 19780
rect 15384 19703 15436 19712
rect 15384 19669 15393 19703
rect 15393 19669 15427 19703
rect 15427 19669 15436 19703
rect 15384 19660 15436 19669
rect 7214 19558 7266 19610
rect 7278 19558 7330 19610
rect 7342 19558 7394 19610
rect 7406 19558 7458 19610
rect 7470 19558 7522 19610
rect 13214 19558 13266 19610
rect 13278 19558 13330 19610
rect 13342 19558 13394 19610
rect 13406 19558 13458 19610
rect 13470 19558 13522 19610
rect 19214 19558 19266 19610
rect 19278 19558 19330 19610
rect 19342 19558 19394 19610
rect 19406 19558 19458 19610
rect 19470 19558 19522 19610
rect 4068 19456 4120 19508
rect 6276 19456 6328 19508
rect 6368 19456 6420 19508
rect 9312 19456 9364 19508
rect 4620 19363 4672 19372
rect 4620 19329 4654 19363
rect 4654 19329 4672 19363
rect 4620 19320 4672 19329
rect 5908 19363 5960 19372
rect 5908 19329 5917 19363
rect 5917 19329 5951 19363
rect 5951 19329 5960 19363
rect 5908 19320 5960 19329
rect 3240 19159 3292 19168
rect 3240 19125 3249 19159
rect 3249 19125 3283 19159
rect 3283 19125 3292 19159
rect 3240 19116 3292 19125
rect 4068 19116 4120 19168
rect 6276 19320 6328 19372
rect 8300 19363 8352 19372
rect 8300 19329 8309 19363
rect 8309 19329 8343 19363
rect 8343 19329 8352 19363
rect 8300 19320 8352 19329
rect 10048 19320 10100 19372
rect 10784 19320 10836 19372
rect 10876 19363 10928 19372
rect 10876 19329 10885 19363
rect 10885 19329 10919 19363
rect 10919 19329 10928 19363
rect 10876 19320 10928 19329
rect 12256 19388 12308 19440
rect 12900 19388 12952 19440
rect 8576 19295 8628 19304
rect 8576 19261 8585 19295
rect 8585 19261 8619 19295
rect 8619 19261 8628 19295
rect 8576 19252 8628 19261
rect 14096 19456 14148 19508
rect 15568 19456 15620 19508
rect 17776 19456 17828 19508
rect 17960 19499 18012 19508
rect 17960 19465 17969 19499
rect 17969 19465 18003 19499
rect 18003 19465 18012 19499
rect 17960 19456 18012 19465
rect 18788 19456 18840 19508
rect 14556 19388 14608 19440
rect 15936 19388 15988 19440
rect 18144 19388 18196 19440
rect 18328 19388 18380 19440
rect 11796 19184 11848 19236
rect 5724 19159 5776 19168
rect 5724 19125 5733 19159
rect 5733 19125 5767 19159
rect 5767 19125 5776 19159
rect 5724 19116 5776 19125
rect 7840 19116 7892 19168
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11152 19159 11204 19168
rect 11152 19125 11161 19159
rect 11161 19125 11195 19159
rect 11195 19125 11204 19159
rect 11152 19116 11204 19125
rect 13820 19116 13872 19168
rect 15016 19320 15068 19372
rect 19616 19388 19668 19440
rect 15200 19184 15252 19236
rect 17960 19116 18012 19168
rect 19800 19116 19852 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 10214 19014 10266 19066
rect 10278 19014 10330 19066
rect 10342 19014 10394 19066
rect 10406 19014 10458 19066
rect 10470 19014 10522 19066
rect 16214 19014 16266 19066
rect 16278 19014 16330 19066
rect 16342 19014 16394 19066
rect 16406 19014 16458 19066
rect 16470 19014 16522 19066
rect 3240 18912 3292 18964
rect 4160 18912 4212 18964
rect 4620 18912 4672 18964
rect 6276 18955 6328 18964
rect 6276 18921 6285 18955
rect 6285 18921 6319 18955
rect 6319 18921 6328 18955
rect 6276 18912 6328 18921
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 8576 18912 8628 18964
rect 10784 18912 10836 18964
rect 5816 18844 5868 18896
rect 7840 18887 7892 18896
rect 7840 18853 7849 18887
rect 7849 18853 7883 18887
rect 7883 18853 7892 18887
rect 7840 18844 7892 18853
rect 5172 18776 5224 18828
rect 5908 18776 5960 18828
rect 9312 18776 9364 18828
rect 12440 18912 12492 18964
rect 12900 18912 12952 18964
rect 13728 18912 13780 18964
rect 5724 18708 5776 18760
rect 5908 18640 5960 18692
rect 11796 18640 11848 18692
rect 14096 18683 14148 18692
rect 14096 18649 14105 18683
rect 14105 18649 14139 18683
rect 14139 18649 14148 18683
rect 14096 18640 14148 18649
rect 14556 18844 14608 18896
rect 16948 18955 17000 18964
rect 16948 18921 16957 18955
rect 16957 18921 16991 18955
rect 16991 18921 17000 18955
rect 16948 18912 17000 18921
rect 18236 18912 18288 18964
rect 19616 18955 19668 18964
rect 19616 18921 19625 18955
rect 19625 18921 19659 18955
rect 19659 18921 19668 18955
rect 19616 18912 19668 18921
rect 15384 18819 15436 18828
rect 15384 18785 15393 18819
rect 15393 18785 15427 18819
rect 15427 18785 15436 18819
rect 15384 18776 15436 18785
rect 15476 18708 15528 18760
rect 16120 18708 16172 18760
rect 2872 18615 2924 18624
rect 2872 18581 2881 18615
rect 2881 18581 2915 18615
rect 2915 18581 2924 18615
rect 2872 18572 2924 18581
rect 14188 18572 14240 18624
rect 14372 18615 14424 18624
rect 14372 18581 14381 18615
rect 14381 18581 14415 18615
rect 14415 18581 14424 18615
rect 14372 18572 14424 18581
rect 14464 18615 14516 18624
rect 14464 18581 14473 18615
rect 14473 18581 14507 18615
rect 14507 18581 14516 18615
rect 14464 18572 14516 18581
rect 17040 18572 17092 18624
rect 18144 18615 18196 18624
rect 18144 18581 18153 18615
rect 18153 18581 18187 18615
rect 18187 18581 18196 18615
rect 18144 18572 18196 18581
rect 19708 18751 19760 18760
rect 19708 18717 19717 18751
rect 19717 18717 19751 18751
rect 19751 18717 19760 18751
rect 19708 18708 19760 18717
rect 19800 18708 19852 18760
rect 19892 18708 19944 18760
rect 7214 18470 7266 18522
rect 7278 18470 7330 18522
rect 7342 18470 7394 18522
rect 7406 18470 7458 18522
rect 7470 18470 7522 18522
rect 13214 18470 13266 18522
rect 13278 18470 13330 18522
rect 13342 18470 13394 18522
rect 13406 18470 13458 18522
rect 13470 18470 13522 18522
rect 19214 18470 19266 18522
rect 19278 18470 19330 18522
rect 19342 18470 19394 18522
rect 19406 18470 19458 18522
rect 19470 18470 19522 18522
rect 4712 18207 4764 18216
rect 4712 18173 4721 18207
rect 4721 18173 4755 18207
rect 4755 18173 4764 18207
rect 4712 18164 4764 18173
rect 9312 18368 9364 18420
rect 8024 18275 8076 18284
rect 8024 18241 8033 18275
rect 8033 18241 8067 18275
rect 8067 18241 8076 18275
rect 8024 18232 8076 18241
rect 10048 18232 10100 18284
rect 12440 18368 12492 18420
rect 14372 18368 14424 18420
rect 14648 18368 14700 18420
rect 14464 18300 14516 18352
rect 14188 18232 14240 18284
rect 15936 18411 15988 18420
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 16948 18368 17000 18420
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 16120 18343 16172 18352
rect 16120 18309 16129 18343
rect 16129 18309 16163 18343
rect 16163 18309 16172 18343
rect 16120 18300 16172 18309
rect 17040 18300 17092 18352
rect 19800 18300 19852 18352
rect 15384 18207 15436 18216
rect 15384 18173 15393 18207
rect 15393 18173 15427 18207
rect 15427 18173 15436 18207
rect 15384 18164 15436 18173
rect 18052 18232 18104 18284
rect 15660 18164 15712 18216
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 14096 18028 14148 18080
rect 14648 18028 14700 18080
rect 16672 18028 16724 18080
rect 16948 18028 17000 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 10214 17926 10266 17978
rect 10278 17926 10330 17978
rect 10342 17926 10394 17978
rect 10406 17926 10458 17978
rect 10470 17926 10522 17978
rect 16214 17926 16266 17978
rect 16278 17926 16330 17978
rect 16342 17926 16394 17978
rect 16406 17926 16458 17978
rect 16470 17926 16522 17978
rect 9312 17824 9364 17876
rect 1860 17688 1912 17740
rect 2136 17688 2188 17740
rect 4712 17688 4764 17740
rect 4804 17688 4856 17740
rect 1584 17663 1636 17672
rect 1584 17629 1593 17663
rect 1593 17629 1627 17663
rect 1627 17629 1636 17663
rect 1584 17620 1636 17629
rect 2964 17527 3016 17536
rect 2964 17493 2973 17527
rect 2973 17493 3007 17527
rect 3007 17493 3016 17527
rect 2964 17484 3016 17493
rect 4068 17484 4120 17536
rect 4804 17552 4856 17604
rect 13728 17824 13780 17876
rect 14188 17867 14240 17876
rect 14188 17833 14197 17867
rect 14197 17833 14231 17867
rect 14231 17833 14240 17867
rect 14188 17824 14240 17833
rect 15384 17824 15436 17876
rect 16120 17824 16172 17876
rect 17960 17824 18012 17876
rect 5816 17663 5868 17672
rect 5816 17629 5825 17663
rect 5825 17629 5859 17663
rect 5859 17629 5868 17663
rect 5816 17620 5868 17629
rect 6552 17552 6604 17604
rect 9312 17620 9364 17672
rect 9772 17552 9824 17604
rect 5816 17484 5868 17536
rect 7564 17527 7616 17536
rect 7564 17493 7573 17527
rect 7573 17493 7607 17527
rect 7607 17493 7616 17527
rect 7564 17484 7616 17493
rect 8668 17527 8720 17536
rect 8668 17493 8677 17527
rect 8677 17493 8711 17527
rect 8711 17493 8720 17527
rect 8668 17484 8720 17493
rect 9404 17484 9456 17536
rect 9496 17527 9548 17536
rect 9496 17493 9505 17527
rect 9505 17493 9539 17527
rect 9539 17493 9548 17527
rect 9496 17484 9548 17493
rect 18052 17688 18104 17740
rect 14372 17620 14424 17672
rect 15660 17620 15712 17672
rect 16948 17663 17000 17672
rect 19800 17688 19852 17740
rect 16948 17629 16966 17663
rect 16966 17629 17000 17663
rect 16948 17620 17000 17629
rect 16672 17552 16724 17604
rect 16856 17552 16908 17604
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 19708 17620 19760 17672
rect 10324 17484 10376 17536
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 11060 17484 11112 17536
rect 19800 17595 19852 17604
rect 19800 17561 19809 17595
rect 19809 17561 19843 17595
rect 19843 17561 19852 17595
rect 19800 17552 19852 17561
rect 18236 17527 18288 17536
rect 18236 17493 18245 17527
rect 18245 17493 18279 17527
rect 18279 17493 18288 17527
rect 18236 17484 18288 17493
rect 7214 17382 7266 17434
rect 7278 17382 7330 17434
rect 7342 17382 7394 17434
rect 7406 17382 7458 17434
rect 7470 17382 7522 17434
rect 13214 17382 13266 17434
rect 13278 17382 13330 17434
rect 13342 17382 13394 17434
rect 13406 17382 13458 17434
rect 13470 17382 13522 17434
rect 19214 17382 19266 17434
rect 19278 17382 19330 17434
rect 19342 17382 19394 17434
rect 19406 17382 19458 17434
rect 19470 17382 19522 17434
rect 5172 17323 5224 17332
rect 5172 17289 5181 17323
rect 5181 17289 5215 17323
rect 5215 17289 5224 17323
rect 5172 17280 5224 17289
rect 6552 17280 6604 17332
rect 8668 17280 8720 17332
rect 1952 17187 2004 17196
rect 1952 17153 1986 17187
rect 1986 17153 2004 17187
rect 1952 17144 2004 17153
rect 3608 17212 3660 17264
rect 10324 17280 10376 17332
rect 12440 17280 12492 17332
rect 15384 17280 15436 17332
rect 16856 17323 16908 17332
rect 16856 17289 16865 17323
rect 16865 17289 16899 17323
rect 16899 17289 16908 17323
rect 18052 17323 18104 17332
rect 16856 17280 16908 17289
rect 18052 17289 18061 17323
rect 18061 17289 18095 17323
rect 18095 17289 18104 17323
rect 18052 17280 18104 17289
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 5172 17144 5224 17196
rect 2964 17076 3016 17128
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 3056 16983 3108 16992
rect 3056 16949 3065 16983
rect 3065 16949 3099 16983
rect 3099 16949 3108 16983
rect 3056 16940 3108 16949
rect 10048 17144 10100 17196
rect 10508 17144 10560 17196
rect 13728 17212 13780 17264
rect 14096 17212 14148 17264
rect 19616 17212 19668 17264
rect 3516 16940 3568 16992
rect 4620 16983 4672 16992
rect 4620 16949 4629 16983
rect 4629 16949 4663 16983
rect 4663 16949 4672 16983
rect 4620 16940 4672 16949
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 7564 17076 7616 17128
rect 8576 17076 8628 17128
rect 9496 17076 9548 17128
rect 11060 17187 11112 17196
rect 11060 17153 11069 17187
rect 11069 17153 11103 17187
rect 11103 17153 11112 17187
rect 11060 17144 11112 17153
rect 12348 17144 12400 17196
rect 7104 16940 7156 16992
rect 8668 16940 8720 16992
rect 10876 16940 10928 16992
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 18328 16983 18380 16992
rect 18328 16949 18337 16983
rect 18337 16949 18371 16983
rect 18371 16949 18380 16983
rect 18328 16940 18380 16949
rect 19800 16940 19852 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 10214 16838 10266 16890
rect 10278 16838 10330 16890
rect 10342 16838 10394 16890
rect 10406 16838 10458 16890
rect 10470 16838 10522 16890
rect 16214 16838 16266 16890
rect 16278 16838 16330 16890
rect 16342 16838 16394 16890
rect 16406 16838 16458 16890
rect 16470 16838 16522 16890
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 3516 16736 3568 16788
rect 3608 16736 3660 16788
rect 3884 16736 3936 16788
rect 4988 16736 5040 16788
rect 10876 16779 10928 16788
rect 2136 16575 2188 16584
rect 2136 16541 2170 16575
rect 2170 16541 2188 16575
rect 2136 16532 2188 16541
rect 3700 16600 3752 16652
rect 3976 16600 4028 16652
rect 10876 16745 10900 16779
rect 10900 16745 10928 16779
rect 10876 16736 10928 16745
rect 12348 16779 12400 16788
rect 12348 16745 12357 16779
rect 12357 16745 12391 16779
rect 12391 16745 12400 16779
rect 12348 16736 12400 16745
rect 13728 16736 13780 16788
rect 8576 16600 8628 16652
rect 10968 16600 11020 16652
rect 15200 16736 15252 16788
rect 16856 16736 16908 16788
rect 17132 16600 17184 16652
rect 3884 16532 3936 16584
rect 5540 16532 5592 16584
rect 14372 16532 14424 16584
rect 15016 16532 15068 16584
rect 15476 16532 15528 16584
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 18328 16532 18380 16584
rect 20260 16532 20312 16584
rect 940 16464 992 16516
rect 1584 16464 1636 16516
rect 3056 16464 3108 16516
rect 3332 16396 3384 16448
rect 3884 16396 3936 16448
rect 3976 16439 4028 16448
rect 3976 16405 4001 16439
rect 4001 16405 4028 16439
rect 4620 16464 4672 16516
rect 3976 16396 4028 16405
rect 7104 16439 7156 16448
rect 7104 16405 7113 16439
rect 7113 16405 7147 16439
rect 7147 16405 7156 16439
rect 7104 16396 7156 16405
rect 7840 16396 7892 16448
rect 13084 16396 13136 16448
rect 14464 16396 14516 16448
rect 15292 16507 15344 16516
rect 15292 16473 15301 16507
rect 15301 16473 15335 16507
rect 15335 16473 15344 16507
rect 15292 16464 15344 16473
rect 16028 16464 16080 16516
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 14832 16439 14884 16448
rect 14832 16405 14841 16439
rect 14841 16405 14875 16439
rect 14875 16405 14884 16439
rect 14832 16396 14884 16405
rect 17868 16396 17920 16448
rect 18972 16439 19024 16448
rect 18972 16405 18981 16439
rect 18981 16405 19015 16439
rect 19015 16405 19024 16439
rect 18972 16396 19024 16405
rect 7214 16294 7266 16346
rect 7278 16294 7330 16346
rect 7342 16294 7394 16346
rect 7406 16294 7458 16346
rect 7470 16294 7522 16346
rect 13214 16294 13266 16346
rect 13278 16294 13330 16346
rect 13342 16294 13394 16346
rect 13406 16294 13458 16346
rect 13470 16294 13522 16346
rect 19214 16294 19266 16346
rect 19278 16294 19330 16346
rect 19342 16294 19394 16346
rect 19406 16294 19458 16346
rect 19470 16294 19522 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 12440 16192 12492 16244
rect 1584 16124 1636 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 10140 16056 10192 16108
rect 10600 16124 10652 16176
rect 14832 16192 14884 16244
rect 15292 16192 15344 16244
rect 15936 16192 15988 16244
rect 12808 16124 12860 16176
rect 14464 16167 14516 16176
rect 14464 16133 14473 16167
rect 14473 16133 14507 16167
rect 14507 16133 14516 16167
rect 14464 16124 14516 16133
rect 14372 16056 14424 16108
rect 16028 16124 16080 16176
rect 18144 16124 18196 16176
rect 18236 16124 18288 16176
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 18972 16056 19024 16108
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 3516 15895 3568 15904
rect 3516 15861 3525 15895
rect 3525 15861 3559 15895
rect 3559 15861 3568 15895
rect 3516 15852 3568 15861
rect 10600 15852 10652 15904
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 14740 15920 14792 15972
rect 17316 15963 17368 15972
rect 17316 15929 17325 15963
rect 17325 15929 17359 15963
rect 17359 15929 17368 15963
rect 18236 16031 18288 16040
rect 18236 15997 18245 16031
rect 18245 15997 18279 16031
rect 18279 15997 18288 16031
rect 18236 15988 18288 15997
rect 17316 15920 17368 15929
rect 15384 15852 15436 15904
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 18696 15895 18748 15904
rect 18696 15861 18705 15895
rect 18705 15861 18739 15895
rect 18739 15861 18748 15895
rect 18696 15852 18748 15861
rect 19616 15852 19668 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 10214 15750 10266 15802
rect 10278 15750 10330 15802
rect 10342 15750 10394 15802
rect 10406 15750 10458 15802
rect 10470 15750 10522 15802
rect 16214 15750 16266 15802
rect 16278 15750 16330 15802
rect 16342 15750 16394 15802
rect 16406 15750 16458 15802
rect 16470 15750 16522 15802
rect 10600 15648 10652 15700
rect 10692 15648 10744 15700
rect 11152 15648 11204 15700
rect 11796 15648 11848 15700
rect 13728 15648 13780 15700
rect 3332 15512 3384 15564
rect 6368 15555 6420 15564
rect 3884 15444 3936 15496
rect 6368 15521 6377 15555
rect 6377 15521 6411 15555
rect 6411 15521 6420 15555
rect 6368 15512 6420 15521
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 1952 15376 2004 15428
rect 3976 15419 4028 15428
rect 3976 15385 3985 15419
rect 3985 15385 4019 15419
rect 4019 15385 4028 15419
rect 3976 15376 4028 15385
rect 3792 15308 3844 15360
rect 4896 15487 4948 15496
rect 4896 15453 4905 15487
rect 4905 15453 4939 15487
rect 4939 15453 4948 15487
rect 4896 15444 4948 15453
rect 11520 15512 11572 15564
rect 14740 15648 14792 15700
rect 15384 15648 15436 15700
rect 15936 15691 15988 15700
rect 15936 15657 15945 15691
rect 15945 15657 15979 15691
rect 15979 15657 15988 15691
rect 15936 15648 15988 15657
rect 17316 15648 17368 15700
rect 17408 15648 17460 15700
rect 18880 15691 18932 15700
rect 18880 15657 18889 15691
rect 18889 15657 18923 15691
rect 18923 15657 18932 15691
rect 18880 15648 18932 15657
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 15476 15623 15528 15632
rect 15476 15589 15485 15623
rect 15485 15589 15519 15623
rect 15519 15589 15528 15623
rect 15476 15580 15528 15589
rect 15660 15623 15712 15632
rect 15660 15589 15669 15623
rect 15669 15589 15703 15623
rect 15703 15589 15712 15623
rect 15660 15580 15712 15589
rect 18328 15580 18380 15632
rect 14096 15555 14148 15564
rect 14096 15521 14105 15555
rect 14105 15521 14139 15555
rect 14139 15521 14148 15555
rect 14096 15512 14148 15521
rect 16028 15555 16080 15564
rect 16028 15521 16037 15555
rect 16037 15521 16071 15555
rect 16071 15521 16080 15555
rect 16028 15512 16080 15521
rect 11060 15444 11112 15496
rect 14832 15444 14884 15496
rect 15568 15444 15620 15496
rect 18236 15444 18288 15496
rect 18696 15444 18748 15496
rect 18788 15487 18840 15496
rect 18788 15453 18797 15487
rect 18797 15453 18831 15487
rect 18831 15453 18840 15487
rect 18788 15444 18840 15453
rect 6184 15376 6236 15428
rect 6644 15419 6696 15428
rect 6644 15385 6653 15419
rect 6653 15385 6687 15419
rect 6687 15385 6696 15419
rect 6644 15376 6696 15385
rect 8024 15376 8076 15428
rect 10232 15376 10284 15428
rect 10692 15376 10744 15428
rect 4712 15351 4764 15360
rect 4712 15317 4721 15351
rect 4721 15317 4755 15351
rect 4755 15317 4764 15351
rect 4712 15308 4764 15317
rect 7656 15308 7708 15360
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 12716 15376 12768 15428
rect 13084 15376 13136 15428
rect 17868 15376 17920 15428
rect 18972 15444 19024 15496
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 11704 15308 11756 15360
rect 16672 15351 16724 15360
rect 16672 15317 16681 15351
rect 16681 15317 16715 15351
rect 16715 15317 16724 15351
rect 16672 15308 16724 15317
rect 18880 15308 18932 15360
rect 19616 15308 19668 15360
rect 7214 15206 7266 15258
rect 7278 15206 7330 15258
rect 7342 15206 7394 15258
rect 7406 15206 7458 15258
rect 7470 15206 7522 15258
rect 13214 15206 13266 15258
rect 13278 15206 13330 15258
rect 13342 15206 13394 15258
rect 13406 15206 13458 15258
rect 13470 15206 13522 15258
rect 19214 15206 19266 15258
rect 19278 15206 19330 15258
rect 19342 15206 19394 15258
rect 19406 15206 19458 15258
rect 19470 15206 19522 15258
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 1952 14900 2004 14952
rect 2320 15079 2372 15088
rect 2320 15045 2329 15079
rect 2329 15045 2363 15079
rect 2363 15045 2372 15079
rect 2320 15036 2372 15045
rect 4896 15104 4948 15156
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 4160 15036 4212 15088
rect 5264 15036 5316 15088
rect 7656 15104 7708 15156
rect 9220 15104 9272 15156
rect 10968 15104 11020 15156
rect 6460 15011 6512 15020
rect 6460 14977 6469 15011
rect 6469 14977 6503 15011
rect 6503 14977 6512 15011
rect 6460 14968 6512 14977
rect 8024 14968 8076 15020
rect 8484 14968 8536 15020
rect 8576 15011 8628 15020
rect 8576 14977 8585 15011
rect 8585 14977 8619 15011
rect 8619 14977 8628 15011
rect 8576 14968 8628 14977
rect 10140 14968 10192 15020
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 3700 14900 3752 14952
rect 3884 14900 3936 14952
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 6184 14943 6236 14952
rect 6184 14909 6193 14943
rect 6193 14909 6227 14943
rect 6227 14909 6236 14943
rect 6184 14900 6236 14909
rect 6736 14943 6788 14952
rect 6736 14909 6745 14943
rect 6745 14909 6779 14943
rect 6779 14909 6788 14943
rect 6736 14900 6788 14909
rect 10232 14900 10284 14952
rect 2136 14764 2188 14816
rect 7748 14764 7800 14816
rect 11152 14943 11204 14952
rect 11152 14909 11160 14943
rect 11160 14909 11194 14943
rect 11194 14909 11204 14943
rect 11152 14900 11204 14909
rect 11796 14900 11848 14952
rect 14096 15147 14148 15156
rect 14096 15113 14105 15147
rect 14105 15113 14139 15147
rect 14139 15113 14148 15147
rect 14096 15104 14148 15113
rect 14372 15147 14424 15156
rect 14372 15113 14381 15147
rect 14381 15113 14415 15147
rect 14415 15113 14424 15147
rect 14372 15104 14424 15113
rect 16672 15104 16724 15156
rect 17132 15147 17184 15156
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 17776 15104 17828 15156
rect 18788 15104 18840 15156
rect 15476 15079 15528 15088
rect 15476 15045 15494 15079
rect 15494 15045 15528 15079
rect 18236 15079 18288 15088
rect 15476 15036 15528 15045
rect 18236 15045 18245 15079
rect 18245 15045 18279 15079
rect 18279 15045 18288 15079
rect 18236 15036 18288 15045
rect 14740 14968 14792 15020
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 18880 14968 18932 15020
rect 20352 15036 20404 15088
rect 18144 14900 18196 14952
rect 17316 14832 17368 14884
rect 17868 14832 17920 14884
rect 12164 14807 12216 14816
rect 12164 14773 12173 14807
rect 12173 14773 12207 14807
rect 12207 14773 12216 14807
rect 12164 14764 12216 14773
rect 12348 14764 12400 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 10214 14662 10266 14714
rect 10278 14662 10330 14714
rect 10342 14662 10394 14714
rect 10406 14662 10458 14714
rect 10470 14662 10522 14714
rect 16214 14662 16266 14714
rect 16278 14662 16330 14714
rect 16342 14662 16394 14714
rect 16406 14662 16458 14714
rect 16470 14662 16522 14714
rect 1492 14560 1544 14612
rect 2320 14560 2372 14612
rect 3700 14560 3752 14612
rect 5264 14560 5316 14612
rect 5908 14560 5960 14612
rect 6460 14560 6512 14612
rect 6736 14603 6788 14612
rect 6736 14569 6745 14603
rect 6745 14569 6779 14603
rect 6779 14569 6788 14603
rect 6736 14560 6788 14569
rect 3792 14467 3844 14476
rect 3792 14433 3801 14467
rect 3801 14433 3835 14467
rect 3835 14433 3844 14467
rect 3792 14424 3844 14433
rect 4712 14424 4764 14476
rect 2780 14356 2832 14408
rect 6276 14424 6328 14476
rect 7748 14560 7800 14612
rect 8576 14560 8628 14612
rect 11336 14560 11388 14612
rect 12164 14560 12216 14612
rect 12256 14560 12308 14612
rect 18604 14560 18656 14612
rect 6368 14356 6420 14408
rect 14740 14535 14792 14544
rect 14740 14501 14749 14535
rect 14749 14501 14783 14535
rect 14783 14501 14792 14535
rect 14740 14492 14792 14501
rect 1952 14288 2004 14340
rect 12256 14424 12308 14476
rect 12348 14424 12400 14476
rect 11336 14356 11388 14408
rect 7012 14220 7064 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 12716 14288 12768 14340
rect 15844 14288 15896 14340
rect 15936 14220 15988 14272
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 7214 14118 7266 14170
rect 7278 14118 7330 14170
rect 7342 14118 7394 14170
rect 7406 14118 7458 14170
rect 7470 14118 7522 14170
rect 13214 14118 13266 14170
rect 13278 14118 13330 14170
rect 13342 14118 13394 14170
rect 13406 14118 13458 14170
rect 13470 14118 13522 14170
rect 19214 14118 19266 14170
rect 19278 14118 19330 14170
rect 19342 14118 19394 14170
rect 19406 14118 19458 14170
rect 19470 14118 19522 14170
rect 2044 14016 2096 14068
rect 7748 14016 7800 14068
rect 8484 14016 8536 14068
rect 6368 13948 6420 14000
rect 6920 13923 6972 13932
rect 6920 13889 6924 13923
rect 6924 13889 6958 13923
rect 6958 13889 6972 13923
rect 6920 13880 6972 13889
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 7840 13948 7892 14000
rect 10692 14016 10744 14068
rect 14096 14059 14148 14068
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 8392 13880 8444 13932
rect 8576 13880 8628 13932
rect 10140 13948 10192 14000
rect 12716 13948 12768 14000
rect 1860 13812 1912 13864
rect 9128 13880 9180 13932
rect 16304 14059 16356 14068
rect 16304 14025 16313 14059
rect 16313 14025 16347 14059
rect 16347 14025 16356 14059
rect 16304 14016 16356 14025
rect 18236 14016 18288 14068
rect 15476 13991 15528 14000
rect 15476 13957 15516 13991
rect 15516 13957 15528 13991
rect 15476 13948 15528 13957
rect 16028 13880 16080 13932
rect 16948 13923 17000 13932
rect 16948 13889 16971 13923
rect 16971 13889 17000 13923
rect 16948 13880 17000 13889
rect 18880 14016 18932 14068
rect 19616 13948 19668 14000
rect 10508 13855 10560 13864
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 15752 13855 15804 13864
rect 15752 13821 15761 13855
rect 15761 13821 15795 13855
rect 15795 13821 15804 13855
rect 15752 13812 15804 13821
rect 15844 13812 15896 13864
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 6736 13719 6788 13728
rect 6736 13685 6745 13719
rect 6745 13685 6779 13719
rect 6779 13685 6788 13719
rect 6736 13676 6788 13685
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 9956 13676 10008 13728
rect 15936 13719 15988 13728
rect 15936 13685 15945 13719
rect 15945 13685 15979 13719
rect 15979 13685 15988 13719
rect 15936 13676 15988 13685
rect 18052 13719 18104 13728
rect 18052 13685 18061 13719
rect 18061 13685 18095 13719
rect 18095 13685 18104 13719
rect 18052 13676 18104 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 10214 13574 10266 13626
rect 10278 13574 10330 13626
rect 10342 13574 10394 13626
rect 10406 13574 10458 13626
rect 10470 13574 10522 13626
rect 16214 13574 16266 13626
rect 16278 13574 16330 13626
rect 16342 13574 16394 13626
rect 16406 13574 16458 13626
rect 16470 13574 16522 13626
rect 6276 13472 6328 13524
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 20260 13472 20312 13524
rect 3148 13447 3200 13456
rect 3148 13413 3157 13447
rect 3157 13413 3191 13447
rect 3191 13413 3200 13447
rect 3148 13404 3200 13413
rect 2044 13336 2096 13388
rect 10692 13404 10744 13456
rect 2780 13268 2832 13320
rect 3332 13268 3384 13320
rect 6920 13336 6972 13388
rect 8760 13336 8812 13388
rect 11428 13336 11480 13388
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 2964 13200 3016 13252
rect 3516 13243 3568 13252
rect 3516 13209 3525 13243
rect 3525 13209 3559 13243
rect 3559 13209 3568 13243
rect 3516 13200 3568 13209
rect 4252 13243 4304 13252
rect 4252 13209 4261 13243
rect 4261 13209 4295 13243
rect 4295 13209 4304 13243
rect 4252 13200 4304 13209
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 15476 13447 15528 13456
rect 15476 13413 15485 13447
rect 15485 13413 15519 13447
rect 15519 13413 15528 13447
rect 15476 13404 15528 13413
rect 16948 13404 17000 13456
rect 14096 13379 14148 13388
rect 14096 13345 14105 13379
rect 14105 13345 14139 13379
rect 14139 13345 14148 13379
rect 14096 13336 14148 13345
rect 15752 13268 15804 13320
rect 15936 13311 15988 13320
rect 15936 13277 15970 13311
rect 15970 13277 15988 13311
rect 15936 13268 15988 13277
rect 16672 13268 16724 13320
rect 19064 13311 19116 13320
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 5724 13200 5776 13252
rect 2320 13132 2372 13184
rect 4528 13132 4580 13184
rect 7012 13200 7064 13252
rect 9128 13200 9180 13252
rect 9496 13200 9548 13252
rect 10508 13200 10560 13252
rect 10876 13200 10928 13252
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9588 13132 9640 13184
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 14740 13200 14792 13252
rect 18328 13200 18380 13252
rect 10692 13132 10744 13141
rect 17408 13132 17460 13184
rect 7214 13030 7266 13082
rect 7278 13030 7330 13082
rect 7342 13030 7394 13082
rect 7406 13030 7458 13082
rect 7470 13030 7522 13082
rect 13214 13030 13266 13082
rect 13278 13030 13330 13082
rect 13342 13030 13394 13082
rect 13406 13030 13458 13082
rect 13470 13030 13522 13082
rect 19214 13030 19266 13082
rect 19278 13030 19330 13082
rect 19342 13030 19394 13082
rect 19406 13030 19458 13082
rect 19470 13030 19522 13082
rect 1676 12928 1728 12980
rect 2320 12928 2372 12980
rect 2504 12724 2556 12776
rect 2964 12860 3016 12912
rect 3332 12860 3384 12912
rect 4528 12928 4580 12980
rect 6644 12928 6696 12980
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 5724 12860 5776 12912
rect 6920 12792 6972 12844
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 8484 12860 8536 12912
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 10876 12928 10928 12980
rect 11152 12860 11204 12912
rect 11428 12928 11480 12980
rect 14740 12971 14792 12980
rect 14740 12937 14749 12971
rect 14749 12937 14783 12971
rect 14783 12937 14792 12971
rect 14740 12928 14792 12937
rect 15476 12928 15528 12980
rect 15844 12971 15896 12980
rect 15844 12937 15853 12971
rect 15853 12937 15887 12971
rect 15887 12937 15896 12971
rect 15844 12928 15896 12937
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 19340 12971 19392 12980
rect 19340 12937 19349 12971
rect 19349 12937 19383 12971
rect 19383 12937 19392 12971
rect 19340 12928 19392 12937
rect 16028 12860 16080 12912
rect 17224 12860 17276 12912
rect 17408 12860 17460 12912
rect 8392 12724 8444 12776
rect 9864 12767 9916 12776
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 9864 12724 9916 12733
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 5724 12656 5776 12708
rect 6460 12656 6512 12708
rect 7012 12656 7064 12708
rect 2136 12588 2188 12640
rect 9956 12588 10008 12640
rect 10508 12588 10560 12640
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 13912 12792 13964 12844
rect 14096 12792 14148 12844
rect 14648 12792 14700 12844
rect 15752 12792 15804 12844
rect 18328 12860 18380 12912
rect 18052 12792 18104 12844
rect 18972 12792 19024 12844
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 16948 12588 17000 12640
rect 17868 12631 17920 12640
rect 17868 12597 17877 12631
rect 17877 12597 17911 12631
rect 17911 12597 17920 12631
rect 17868 12588 17920 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 10214 12486 10266 12538
rect 10278 12486 10330 12538
rect 10342 12486 10394 12538
rect 10406 12486 10458 12538
rect 10470 12486 10522 12538
rect 16214 12486 16266 12538
rect 16278 12486 16330 12538
rect 16342 12486 16394 12538
rect 16406 12486 16458 12538
rect 16470 12486 16522 12538
rect 2872 12384 2924 12436
rect 4068 12384 4120 12436
rect 4712 12427 4764 12436
rect 4712 12393 4721 12427
rect 4721 12393 4755 12427
rect 4755 12393 4764 12427
rect 4712 12384 4764 12393
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 9864 12384 9916 12436
rect 10876 12384 10928 12436
rect 11520 12384 11572 12436
rect 3148 12248 3200 12300
rect 3884 12316 3936 12368
rect 1860 12223 1912 12232
rect 1860 12189 1869 12223
rect 1869 12189 1903 12223
rect 1903 12189 1912 12223
rect 1860 12180 1912 12189
rect 3240 12180 3292 12232
rect 2136 12112 2188 12164
rect 4528 12223 4580 12232
rect 4528 12189 4537 12223
rect 4537 12189 4571 12223
rect 4571 12189 4580 12223
rect 10784 12248 10836 12300
rect 4528 12180 4580 12189
rect 9496 12180 9548 12232
rect 10692 12180 10744 12232
rect 13360 12384 13412 12436
rect 13912 12384 13964 12436
rect 11244 12180 11296 12232
rect 12440 12223 12492 12232
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 12440 12180 12492 12189
rect 14096 12359 14148 12368
rect 14096 12325 14105 12359
rect 14105 12325 14139 12359
rect 14139 12325 14148 12359
rect 14096 12316 14148 12325
rect 14740 12316 14792 12368
rect 15200 12316 15252 12368
rect 18328 12384 18380 12436
rect 18880 12427 18932 12436
rect 18880 12393 18889 12427
rect 18889 12393 18923 12427
rect 18923 12393 18932 12427
rect 18880 12384 18932 12393
rect 16948 12291 17000 12300
rect 16948 12257 16957 12291
rect 16957 12257 16991 12291
rect 16991 12257 17000 12291
rect 16948 12248 17000 12257
rect 19340 12248 19392 12300
rect 15568 12180 15620 12232
rect 15844 12155 15896 12164
rect 15844 12121 15853 12155
rect 15853 12121 15887 12155
rect 15887 12121 15896 12155
rect 15844 12112 15896 12121
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 16396 12223 16448 12232
rect 16396 12189 16405 12223
rect 16405 12189 16439 12223
rect 16439 12189 16448 12223
rect 16396 12180 16448 12189
rect 17224 12223 17276 12232
rect 17224 12189 17258 12223
rect 17258 12189 17276 12223
rect 17224 12180 17276 12189
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 19616 12180 19668 12232
rect 5448 12044 5500 12096
rect 8760 12044 8812 12096
rect 12532 12044 12584 12096
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 18328 12087 18380 12096
rect 18328 12053 18337 12087
rect 18337 12053 18371 12087
rect 18371 12053 18380 12087
rect 18328 12044 18380 12053
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 7214 11942 7266 11994
rect 7278 11942 7330 11994
rect 7342 11942 7394 11994
rect 7406 11942 7458 11994
rect 7470 11942 7522 11994
rect 13214 11942 13266 11994
rect 13278 11942 13330 11994
rect 13342 11942 13394 11994
rect 13406 11942 13458 11994
rect 13470 11942 13522 11994
rect 19214 11942 19266 11994
rect 19278 11942 19330 11994
rect 19342 11942 19394 11994
rect 19406 11942 19458 11994
rect 19470 11942 19522 11994
rect 2136 11840 2188 11892
rect 2504 11883 2556 11892
rect 2504 11849 2513 11883
rect 2513 11849 2547 11883
rect 2547 11849 2556 11883
rect 2504 11840 2556 11849
rect 4528 11840 4580 11892
rect 15200 11840 15252 11892
rect 15568 11840 15620 11892
rect 13820 11815 13872 11824
rect 13820 11781 13829 11815
rect 13829 11781 13863 11815
rect 13863 11781 13872 11815
rect 13820 11772 13872 11781
rect 14464 11772 14516 11824
rect 15292 11772 15344 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 12532 11704 12584 11756
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 15844 11883 15896 11892
rect 15844 11849 15853 11883
rect 15853 11849 15887 11883
rect 15887 11849 15896 11883
rect 15844 11840 15896 11849
rect 16212 11840 16264 11892
rect 16396 11840 16448 11892
rect 16672 11840 16724 11892
rect 16948 11815 17000 11824
rect 16948 11781 16957 11815
rect 16957 11781 16991 11815
rect 16991 11781 17000 11815
rect 16948 11772 17000 11781
rect 17316 11815 17368 11824
rect 17316 11781 17325 11815
rect 17325 11781 17359 11815
rect 17359 11781 17368 11815
rect 17316 11772 17368 11781
rect 18512 11840 18564 11892
rect 18880 11883 18932 11892
rect 18880 11849 18889 11883
rect 18889 11849 18923 11883
rect 18923 11849 18932 11883
rect 18880 11840 18932 11849
rect 19064 11840 19116 11892
rect 20076 11840 20128 11892
rect 17776 11679 17828 11688
rect 17776 11645 17785 11679
rect 17785 11645 17819 11679
rect 17819 11645 17828 11679
rect 17776 11636 17828 11645
rect 19616 11772 19668 11824
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 13912 11543 13964 11552
rect 13912 11509 13921 11543
rect 13921 11509 13955 11543
rect 13955 11509 13964 11543
rect 13912 11500 13964 11509
rect 16120 11543 16172 11552
rect 16120 11509 16129 11543
rect 16129 11509 16163 11543
rect 16163 11509 16172 11543
rect 16120 11500 16172 11509
rect 18880 11636 18932 11688
rect 18328 11500 18380 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 10214 11398 10266 11450
rect 10278 11398 10330 11450
rect 10342 11398 10394 11450
rect 10406 11398 10458 11450
rect 10470 11398 10522 11450
rect 16214 11398 16266 11450
rect 16278 11398 16330 11450
rect 16342 11398 16394 11450
rect 16406 11398 16458 11450
rect 16470 11398 16522 11450
rect 3240 11228 3292 11280
rect 2780 11160 2832 11212
rect 5448 11160 5500 11212
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 9220 11296 9272 11348
rect 9588 11339 9640 11348
rect 9588 11305 9597 11339
rect 9597 11305 9631 11339
rect 9631 11305 9640 11339
rect 9588 11296 9640 11305
rect 11060 11296 11112 11348
rect 11520 11296 11572 11348
rect 12440 11296 12492 11348
rect 12532 11339 12584 11348
rect 12532 11305 12541 11339
rect 12541 11305 12575 11339
rect 12575 11305 12584 11339
rect 12532 11296 12584 11305
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 10048 11160 10100 11212
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 3976 11067 4028 11076
rect 3976 11033 3985 11067
rect 3985 11033 4019 11067
rect 4019 11033 4028 11067
rect 3976 11024 4028 11033
rect 4620 11024 4672 11076
rect 4712 11067 4764 11076
rect 4712 11033 4721 11067
rect 4721 11033 4755 11067
rect 4755 11033 4764 11067
rect 4712 11024 4764 11033
rect 8392 11024 8444 11076
rect 8668 11024 8720 11076
rect 9864 11067 9916 11076
rect 9864 11033 9873 11067
rect 9873 11033 9907 11067
rect 9907 11033 9916 11067
rect 9864 11024 9916 11033
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 16948 11160 17000 11212
rect 13820 11092 13872 11144
rect 14648 11092 14700 11144
rect 2320 10956 2372 11008
rect 2688 10999 2740 11008
rect 2688 10965 2697 10999
rect 2697 10965 2731 10999
rect 2731 10965 2740 10999
rect 2688 10956 2740 10965
rect 4528 10956 4580 11008
rect 5356 10956 5408 11008
rect 5724 10956 5776 11008
rect 8300 10999 8352 11008
rect 8300 10965 8309 10999
rect 8309 10965 8343 10999
rect 8343 10965 8352 10999
rect 8300 10956 8352 10965
rect 9036 10956 9088 11008
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 16120 11024 16172 11076
rect 16304 11024 16356 11076
rect 15016 10999 15068 11008
rect 15016 10965 15025 10999
rect 15025 10965 15059 10999
rect 15059 10965 15068 10999
rect 15016 10956 15068 10965
rect 15292 10999 15344 11008
rect 15292 10965 15301 10999
rect 15301 10965 15335 10999
rect 15335 10965 15344 10999
rect 15292 10956 15344 10965
rect 7214 10854 7266 10906
rect 7278 10854 7330 10906
rect 7342 10854 7394 10906
rect 7406 10854 7458 10906
rect 7470 10854 7522 10906
rect 13214 10854 13266 10906
rect 13278 10854 13330 10906
rect 13342 10854 13394 10906
rect 13406 10854 13458 10906
rect 13470 10854 13522 10906
rect 19214 10854 19266 10906
rect 19278 10854 19330 10906
rect 19342 10854 19394 10906
rect 19406 10854 19458 10906
rect 19470 10854 19522 10906
rect 2320 10752 2372 10804
rect 3976 10752 4028 10804
rect 4712 10752 4764 10804
rect 5264 10752 5316 10804
rect 2504 10684 2556 10736
rect 3240 10684 3292 10736
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 5724 10727 5776 10736
rect 5724 10693 5733 10727
rect 5733 10693 5767 10727
rect 5767 10693 5776 10727
rect 5724 10684 5776 10693
rect 9220 10752 9272 10804
rect 9864 10795 9916 10804
rect 9864 10761 9873 10795
rect 9873 10761 9907 10795
rect 9907 10761 9916 10795
rect 9864 10752 9916 10761
rect 10876 10752 10928 10804
rect 11152 10795 11204 10804
rect 11152 10761 11161 10795
rect 11161 10761 11195 10795
rect 11195 10761 11204 10795
rect 11152 10752 11204 10761
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 4068 10412 4120 10464
rect 4804 10591 4856 10600
rect 4804 10557 4813 10591
rect 4813 10557 4847 10591
rect 4847 10557 4856 10591
rect 4804 10548 4856 10557
rect 4620 10480 4672 10532
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 9036 10684 9088 10736
rect 12164 10752 12216 10804
rect 12716 10752 12768 10804
rect 11336 10684 11388 10736
rect 6920 10548 6972 10600
rect 7748 10616 7800 10668
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 13820 10752 13872 10804
rect 16304 10795 16356 10804
rect 16304 10761 16313 10795
rect 16313 10761 16347 10795
rect 16347 10761 16356 10795
rect 16304 10752 16356 10761
rect 16948 10795 17000 10804
rect 16948 10761 16957 10795
rect 16957 10761 16991 10795
rect 16991 10761 17000 10795
rect 16948 10752 17000 10761
rect 15292 10684 15344 10736
rect 15016 10616 15068 10668
rect 15476 10616 15528 10668
rect 18512 10684 18564 10736
rect 18236 10616 18288 10668
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 8300 10548 8352 10600
rect 10048 10548 10100 10600
rect 10140 10548 10192 10600
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 10968 10548 11020 10600
rect 4712 10412 4764 10464
rect 5448 10412 5500 10464
rect 6736 10412 6788 10464
rect 7380 10412 7432 10464
rect 18328 10412 18380 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 10214 10310 10266 10362
rect 10278 10310 10330 10362
rect 10342 10310 10394 10362
rect 10406 10310 10458 10362
rect 10470 10310 10522 10362
rect 16214 10310 16266 10362
rect 16278 10310 16330 10362
rect 16342 10310 16394 10362
rect 16406 10310 16458 10362
rect 16470 10310 16522 10362
rect 1584 10208 1636 10260
rect 2688 10208 2740 10260
rect 2872 10208 2924 10260
rect 3976 10208 4028 10260
rect 4804 10208 4856 10260
rect 5264 10208 5316 10260
rect 5448 10208 5500 10260
rect 5724 10208 5776 10260
rect 2504 10072 2556 10124
rect 3240 10004 3292 10056
rect 4620 10072 4672 10124
rect 4804 10072 4856 10124
rect 4712 9979 4764 9988
rect 1676 9911 1728 9920
rect 1676 9877 1685 9911
rect 1685 9877 1719 9911
rect 1719 9877 1728 9911
rect 1676 9868 1728 9877
rect 4712 9945 4721 9979
rect 4721 9945 4755 9979
rect 4755 9945 4764 9979
rect 4712 9936 4764 9945
rect 5356 10072 5408 10124
rect 5724 10115 5776 10124
rect 5724 10081 5733 10115
rect 5733 10081 5767 10115
rect 5767 10081 5776 10115
rect 5724 10072 5776 10081
rect 6368 10140 6420 10192
rect 6644 10140 6696 10192
rect 8484 10208 8536 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 15476 10251 15528 10260
rect 15476 10217 15485 10251
rect 15485 10217 15519 10251
rect 15519 10217 15528 10251
rect 15476 10208 15528 10217
rect 7380 10072 7432 10124
rect 9772 10072 9824 10124
rect 11520 10072 11572 10124
rect 12440 10072 12492 10124
rect 16948 10208 17000 10260
rect 18144 10208 18196 10260
rect 18052 10072 18104 10124
rect 18696 10115 18748 10124
rect 18696 10081 18705 10115
rect 18705 10081 18739 10115
rect 18739 10081 18748 10115
rect 18696 10072 18748 10081
rect 20444 10115 20496 10124
rect 20444 10081 20453 10115
rect 20453 10081 20487 10115
rect 20487 10081 20496 10115
rect 20444 10072 20496 10081
rect 5264 9936 5316 9988
rect 6092 9936 6144 9988
rect 6460 9936 6512 9988
rect 7748 9936 7800 9988
rect 8208 10004 8260 10056
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 9496 10004 9548 10056
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 10324 10004 10376 10056
rect 12164 10004 12216 10056
rect 18328 10004 18380 10056
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 4068 9868 4120 9920
rect 5080 9868 5132 9920
rect 9312 9868 9364 9920
rect 10048 9868 10100 9920
rect 11612 9979 11664 9988
rect 11612 9945 11621 9979
rect 11621 9945 11655 9979
rect 11655 9945 11664 9979
rect 11612 9936 11664 9945
rect 14372 9979 14424 9988
rect 14372 9945 14406 9979
rect 14406 9945 14424 9979
rect 14372 9936 14424 9945
rect 18880 9979 18932 9988
rect 18880 9945 18889 9979
rect 18889 9945 18923 9979
rect 18923 9945 18932 9979
rect 18880 9936 18932 9945
rect 17960 9911 18012 9920
rect 17960 9877 17969 9911
rect 17969 9877 18003 9911
rect 18003 9877 18012 9911
rect 17960 9868 18012 9877
rect 7214 9766 7266 9818
rect 7278 9766 7330 9818
rect 7342 9766 7394 9818
rect 7406 9766 7458 9818
rect 7470 9766 7522 9818
rect 13214 9766 13266 9818
rect 13278 9766 13330 9818
rect 13342 9766 13394 9818
rect 13406 9766 13458 9818
rect 13470 9766 13522 9818
rect 19214 9766 19266 9818
rect 19278 9766 19330 9818
rect 19342 9766 19394 9818
rect 19406 9766 19458 9818
rect 19470 9766 19522 9818
rect 2504 9707 2556 9716
rect 2504 9673 2513 9707
rect 2513 9673 2547 9707
rect 2547 9673 2556 9707
rect 2504 9664 2556 9673
rect 6552 9664 6604 9716
rect 7748 9707 7800 9716
rect 7748 9673 7757 9707
rect 7757 9673 7791 9707
rect 7791 9673 7800 9707
rect 7748 9664 7800 9673
rect 3792 9639 3844 9648
rect 3792 9605 3801 9639
rect 3801 9605 3835 9639
rect 3835 9605 3844 9639
rect 3792 9596 3844 9605
rect 5540 9596 5592 9648
rect 6276 9596 6328 9648
rect 1676 9528 1728 9580
rect 6092 9528 6144 9580
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 5080 9392 5132 9444
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7748 9528 7800 9580
rect 8208 9596 8260 9648
rect 9772 9664 9824 9716
rect 10324 9707 10376 9716
rect 10324 9673 10333 9707
rect 10333 9673 10367 9707
rect 10367 9673 10376 9707
rect 10324 9664 10376 9673
rect 15016 9664 15068 9716
rect 18420 9664 18472 9716
rect 7932 9571 7984 9580
rect 7932 9537 7941 9571
rect 7941 9537 7975 9571
rect 7975 9537 7984 9571
rect 7932 9528 7984 9537
rect 8116 9528 8168 9580
rect 14372 9596 14424 9648
rect 18880 9596 18932 9648
rect 9956 9528 10008 9580
rect 14188 9528 14240 9580
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 17960 9528 18012 9580
rect 18328 9528 18380 9580
rect 20076 9528 20128 9580
rect 8300 9460 8352 9512
rect 8484 9460 8536 9512
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 18880 9460 18932 9512
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 4804 9324 4856 9376
rect 6644 9324 6696 9376
rect 18788 9392 18840 9444
rect 8576 9324 8628 9376
rect 9864 9324 9916 9376
rect 18512 9324 18564 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 10214 9222 10266 9274
rect 10278 9222 10330 9274
rect 10342 9222 10394 9274
rect 10406 9222 10458 9274
rect 10470 9222 10522 9274
rect 16214 9222 16266 9274
rect 16278 9222 16330 9274
rect 16342 9222 16394 9274
rect 16406 9222 16458 9274
rect 16470 9222 16522 9274
rect 2228 9120 2280 9172
rect 3332 9120 3384 9172
rect 6184 9120 6236 9172
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 8300 9120 8352 9172
rect 17408 9163 17460 9172
rect 17408 9129 17417 9163
rect 17417 9129 17451 9163
rect 17451 9129 17460 9163
rect 17408 9120 17460 9129
rect 17960 9120 18012 9172
rect 18696 9120 18748 9172
rect 20076 9120 20128 9172
rect 6920 9052 6972 9104
rect 8484 9052 8536 9104
rect 4436 8984 4488 9036
rect 5080 8984 5132 9036
rect 5264 8984 5316 9036
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 6368 8916 6420 8968
rect 7748 8984 7800 9036
rect 17868 9052 17920 9104
rect 18972 9052 19024 9104
rect 6736 8848 6788 8900
rect 7564 8916 7616 8968
rect 7932 8916 7984 8968
rect 18512 8984 18564 9036
rect 9680 8916 9732 8968
rect 14096 8959 14148 8968
rect 1676 8823 1728 8832
rect 1676 8789 1685 8823
rect 1685 8789 1719 8823
rect 1719 8789 1728 8823
rect 1676 8780 1728 8789
rect 4344 8780 4396 8832
rect 4988 8780 5040 8832
rect 7012 8780 7064 8832
rect 7104 8780 7156 8832
rect 7656 8780 7708 8832
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 8116 8780 8168 8832
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 14372 8959 14424 8968
rect 14372 8925 14406 8959
rect 14406 8925 14424 8959
rect 14372 8916 14424 8925
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 10784 8848 10836 8900
rect 13728 8848 13780 8900
rect 16856 8891 16908 8900
rect 16856 8857 16874 8891
rect 16874 8857 16908 8891
rect 16856 8848 16908 8857
rect 11060 8780 11112 8832
rect 12164 8780 12216 8832
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 18512 8891 18564 8900
rect 18512 8857 18521 8891
rect 18521 8857 18555 8891
rect 18555 8857 18564 8891
rect 18512 8848 18564 8857
rect 20352 8848 20404 8900
rect 18788 8823 18840 8832
rect 18788 8789 18797 8823
rect 18797 8789 18831 8823
rect 18831 8789 18840 8823
rect 18788 8780 18840 8789
rect 18880 8823 18932 8832
rect 18880 8789 18889 8823
rect 18889 8789 18923 8823
rect 18923 8789 18932 8823
rect 18880 8780 18932 8789
rect 7214 8678 7266 8730
rect 7278 8678 7330 8730
rect 7342 8678 7394 8730
rect 7406 8678 7458 8730
rect 7470 8678 7522 8730
rect 13214 8678 13266 8730
rect 13278 8678 13330 8730
rect 13342 8678 13394 8730
rect 13406 8678 13458 8730
rect 13470 8678 13522 8730
rect 19214 8678 19266 8730
rect 19278 8678 19330 8730
rect 19342 8678 19394 8730
rect 19406 8678 19458 8730
rect 19470 8678 19522 8730
rect 3792 8576 3844 8628
rect 4344 8576 4396 8628
rect 4436 8576 4488 8628
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 4804 8576 4856 8628
rect 4988 8551 5040 8560
rect 4988 8517 4997 8551
rect 4997 8517 5031 8551
rect 5031 8517 5040 8551
rect 4988 8508 5040 8517
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 4160 8372 4212 8424
rect 5264 8576 5316 8628
rect 5724 8576 5776 8628
rect 6184 8576 6236 8628
rect 7472 8508 7524 8560
rect 9312 8551 9364 8560
rect 9312 8517 9321 8551
rect 9321 8517 9355 8551
rect 9355 8517 9364 8551
rect 9312 8508 9364 8517
rect 6184 8440 6236 8492
rect 6276 8440 6328 8492
rect 10784 8576 10836 8628
rect 11060 8576 11112 8628
rect 11244 8619 11296 8628
rect 11244 8585 11261 8619
rect 11261 8585 11295 8619
rect 11295 8585 11296 8619
rect 11244 8576 11296 8585
rect 12440 8576 12492 8628
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 5908 8372 5960 8381
rect 7288 8372 7340 8424
rect 8484 8372 8536 8424
rect 2412 8279 2464 8288
rect 2412 8245 2421 8279
rect 2421 8245 2455 8279
rect 2455 8245 2464 8279
rect 2412 8236 2464 8245
rect 3884 8279 3936 8288
rect 3884 8245 3893 8279
rect 3893 8245 3927 8279
rect 3927 8245 3936 8279
rect 3884 8236 3936 8245
rect 5172 8236 5224 8288
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 5540 8236 5592 8245
rect 7748 8304 7800 8356
rect 8300 8304 8352 8356
rect 9680 8347 9732 8356
rect 9680 8313 9689 8347
rect 9689 8313 9723 8347
rect 9723 8313 9732 8347
rect 9680 8304 9732 8313
rect 10784 8440 10836 8492
rect 11612 8440 11664 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 13728 8440 13780 8492
rect 15476 8508 15528 8560
rect 15752 8508 15804 8560
rect 13820 8415 13872 8424
rect 13820 8381 13829 8415
rect 13829 8381 13863 8415
rect 13863 8381 13872 8415
rect 13820 8372 13872 8381
rect 17592 8576 17644 8628
rect 19248 8508 19300 8560
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 18144 8483 18196 8492
rect 18144 8449 18178 8483
rect 18178 8449 18196 8483
rect 18144 8440 18196 8449
rect 18880 8440 18932 8492
rect 5816 8279 5868 8288
rect 5816 8245 5825 8279
rect 5825 8245 5859 8279
rect 5859 8245 5868 8279
rect 5816 8236 5868 8245
rect 7196 8236 7248 8288
rect 7840 8236 7892 8288
rect 8944 8236 8996 8288
rect 9588 8236 9640 8288
rect 11336 8236 11388 8288
rect 16856 8279 16908 8288
rect 16856 8245 16865 8279
rect 16865 8245 16899 8279
rect 16899 8245 16908 8279
rect 16856 8236 16908 8245
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 18052 8236 18104 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 10214 8134 10266 8186
rect 10278 8134 10330 8186
rect 10342 8134 10394 8186
rect 10406 8134 10458 8186
rect 10470 8134 10522 8186
rect 16214 8134 16266 8186
rect 16278 8134 16330 8186
rect 16342 8134 16394 8186
rect 16406 8134 16458 8186
rect 16470 8134 16522 8186
rect 3884 8032 3936 8084
rect 5356 8032 5408 8084
rect 5816 8032 5868 8084
rect 6736 8032 6788 8084
rect 7288 8075 7340 8084
rect 7288 8041 7297 8075
rect 7297 8041 7331 8075
rect 7331 8041 7340 8075
rect 7288 8032 7340 8041
rect 7564 8075 7616 8084
rect 7564 8041 7573 8075
rect 7573 8041 7607 8075
rect 7607 8041 7616 8075
rect 7564 8032 7616 8041
rect 7656 8032 7708 8084
rect 7840 8032 7892 8084
rect 8208 8075 8260 8084
rect 8208 8041 8217 8075
rect 8217 8041 8251 8075
rect 8251 8041 8260 8075
rect 8208 8032 8260 8041
rect 2228 7896 2280 7948
rect 2504 7896 2556 7948
rect 3148 7896 3200 7948
rect 3148 7692 3200 7744
rect 3700 7760 3752 7812
rect 4804 7896 4856 7948
rect 5540 7896 5592 7948
rect 6184 7964 6236 8016
rect 6736 7896 6788 7948
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6000 7828 6052 7837
rect 6092 7828 6144 7880
rect 4068 7803 4120 7812
rect 4068 7769 4077 7803
rect 4077 7769 4111 7803
rect 4111 7769 4120 7803
rect 4068 7760 4120 7769
rect 4804 7760 4856 7812
rect 5908 7803 5960 7812
rect 5908 7769 5917 7803
rect 5917 7769 5951 7803
rect 5951 7769 5960 7803
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 7196 7828 7248 7880
rect 7564 7896 7616 7948
rect 9680 7896 9732 7948
rect 11704 8032 11756 8084
rect 13820 8032 13872 8084
rect 16856 8032 16908 8084
rect 18144 8032 18196 8084
rect 11336 8007 11388 8016
rect 11336 7973 11345 8007
rect 11345 7973 11379 8007
rect 11379 7973 11388 8007
rect 11336 7964 11388 7973
rect 17868 7964 17920 8016
rect 19248 8075 19300 8084
rect 19248 8041 19257 8075
rect 19257 8041 19291 8075
rect 19291 8041 19300 8075
rect 19248 8032 19300 8041
rect 12164 7896 12216 7948
rect 12440 7896 12492 7948
rect 5908 7760 5960 7769
rect 3976 7692 4028 7744
rect 6184 7735 6236 7744
rect 6184 7701 6193 7735
rect 6193 7701 6227 7735
rect 6227 7701 6236 7735
rect 6184 7692 6236 7701
rect 6644 7760 6696 7812
rect 6920 7803 6972 7812
rect 6920 7769 6929 7803
rect 6929 7769 6963 7803
rect 6963 7769 6972 7803
rect 6920 7760 6972 7769
rect 7012 7692 7064 7744
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 19524 7896 19576 7948
rect 19708 7896 19760 7948
rect 14096 7828 14148 7880
rect 7932 7760 7984 7812
rect 8484 7760 8536 7812
rect 9404 7760 9456 7812
rect 9588 7692 9640 7744
rect 11060 7803 11112 7812
rect 11060 7769 11069 7803
rect 11069 7769 11103 7803
rect 11103 7769 11112 7803
rect 11060 7760 11112 7769
rect 13728 7760 13780 7812
rect 15476 7828 15528 7880
rect 18972 7828 19024 7880
rect 19616 7828 19668 7880
rect 18604 7760 18656 7812
rect 15016 7692 15068 7744
rect 19524 7735 19576 7744
rect 19524 7701 19533 7735
rect 19533 7701 19567 7735
rect 19567 7701 19576 7735
rect 19524 7692 19576 7701
rect 20352 8075 20404 8084
rect 20352 8041 20361 8075
rect 20361 8041 20395 8075
rect 20395 8041 20404 8075
rect 20352 8032 20404 8041
rect 7214 7590 7266 7642
rect 7278 7590 7330 7642
rect 7342 7590 7394 7642
rect 7406 7590 7458 7642
rect 7470 7590 7522 7642
rect 13214 7590 13266 7642
rect 13278 7590 13330 7642
rect 13342 7590 13394 7642
rect 13406 7590 13458 7642
rect 13470 7590 13522 7642
rect 19214 7590 19266 7642
rect 19278 7590 19330 7642
rect 19342 7590 19394 7642
rect 19406 7590 19458 7642
rect 19470 7590 19522 7642
rect 3700 7531 3752 7540
rect 3700 7497 3709 7531
rect 3709 7497 3743 7531
rect 3743 7497 3752 7531
rect 3700 7488 3752 7497
rect 4068 7488 4120 7540
rect 2412 7463 2464 7472
rect 2412 7429 2421 7463
rect 2421 7429 2455 7463
rect 2455 7429 2464 7463
rect 2412 7420 2464 7429
rect 6000 7488 6052 7540
rect 6184 7488 6236 7540
rect 6920 7488 6972 7540
rect 8576 7531 8628 7540
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 11796 7488 11848 7540
rect 18604 7531 18656 7540
rect 18604 7497 18613 7531
rect 18613 7497 18647 7531
rect 18647 7497 18656 7531
rect 18604 7488 18656 7497
rect 18972 7488 19024 7540
rect 7104 7420 7156 7472
rect 1584 7327 1636 7336
rect 1584 7293 1593 7327
rect 1593 7293 1627 7327
rect 1627 7293 1636 7327
rect 1584 7284 1636 7293
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 5540 7352 5592 7404
rect 6276 7352 6328 7404
rect 8944 7352 8996 7404
rect 9588 7420 9640 7472
rect 10140 7463 10192 7472
rect 10140 7429 10149 7463
rect 10149 7429 10183 7463
rect 10183 7429 10192 7463
rect 10140 7420 10192 7429
rect 15752 7420 15804 7472
rect 18420 7463 18472 7472
rect 18420 7429 18429 7463
rect 18429 7429 18463 7463
rect 18463 7429 18472 7463
rect 18420 7420 18472 7429
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 9680 7352 9732 7404
rect 11612 7352 11664 7404
rect 15016 7352 15068 7404
rect 19708 7395 19760 7404
rect 19708 7361 19726 7395
rect 19726 7361 19760 7395
rect 19708 7352 19760 7361
rect 6092 7284 6144 7336
rect 6644 7148 6696 7200
rect 7012 7148 7064 7200
rect 9404 7148 9456 7200
rect 13728 7148 13780 7200
rect 16120 7148 16172 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 10214 7046 10266 7098
rect 10278 7046 10330 7098
rect 10342 7046 10394 7098
rect 10406 7046 10458 7098
rect 10470 7046 10522 7098
rect 16214 7046 16266 7098
rect 16278 7046 16330 7098
rect 16342 7046 16394 7098
rect 16406 7046 16458 7098
rect 16470 7046 16522 7098
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 17408 6944 17460 6996
rect 17684 6987 17736 6996
rect 17684 6953 17693 6987
rect 17693 6953 17727 6987
rect 17727 6953 17736 6987
rect 17684 6944 17736 6953
rect 18420 6987 18472 6996
rect 18420 6953 18429 6987
rect 18429 6953 18463 6987
rect 18463 6953 18472 6987
rect 18420 6944 18472 6953
rect 15016 6876 15068 6928
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 16672 6808 16724 6860
rect 1492 6715 1544 6724
rect 1492 6681 1501 6715
rect 1501 6681 1535 6715
rect 1535 6681 1544 6715
rect 1492 6672 1544 6681
rect 16120 6740 16172 6792
rect 16948 6740 17000 6792
rect 16580 6672 16632 6724
rect 18144 6740 18196 6792
rect 17316 6715 17368 6724
rect 17316 6681 17325 6715
rect 17325 6681 17359 6715
rect 17359 6681 17368 6715
rect 17316 6672 17368 6681
rect 17960 6672 18012 6724
rect 12900 6647 12952 6656
rect 12900 6613 12909 6647
rect 12909 6613 12943 6647
rect 12943 6613 12952 6647
rect 12900 6604 12952 6613
rect 17040 6604 17092 6656
rect 17684 6604 17736 6656
rect 7214 6502 7266 6554
rect 7278 6502 7330 6554
rect 7342 6502 7394 6554
rect 7406 6502 7458 6554
rect 7470 6502 7522 6554
rect 13214 6502 13266 6554
rect 13278 6502 13330 6554
rect 13342 6502 13394 6554
rect 13406 6502 13458 6554
rect 13470 6502 13522 6554
rect 19214 6502 19266 6554
rect 19278 6502 19330 6554
rect 19342 6502 19394 6554
rect 19406 6502 19458 6554
rect 19470 6502 19522 6554
rect 6276 6400 6328 6452
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 9588 6400 9640 6452
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 2872 6264 2924 6316
rect 3976 6264 4028 6316
rect 6920 6264 6972 6316
rect 7564 6264 7616 6316
rect 12808 6400 12860 6452
rect 12900 6400 12952 6452
rect 13728 6264 13780 6316
rect 17040 6400 17092 6452
rect 17684 6400 17736 6452
rect 18144 6400 18196 6452
rect 8024 6239 8076 6248
rect 8024 6205 8033 6239
rect 8033 6205 8067 6239
rect 8067 6205 8076 6239
rect 8024 6196 8076 6205
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 12624 6239 12676 6248
rect 12624 6205 12633 6239
rect 12633 6205 12667 6239
rect 12667 6205 12676 6239
rect 12624 6196 12676 6205
rect 2596 6103 2648 6112
rect 2596 6069 2605 6103
rect 2605 6069 2639 6103
rect 2639 6069 2648 6103
rect 2596 6060 2648 6069
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 10692 6103 10744 6112
rect 10692 6069 10701 6103
rect 10701 6069 10735 6103
rect 10735 6069 10744 6103
rect 10692 6060 10744 6069
rect 12992 6060 13044 6112
rect 16580 6060 16632 6112
rect 18144 6060 18196 6112
rect 18328 6264 18380 6316
rect 19616 6103 19668 6112
rect 19616 6069 19625 6103
rect 19625 6069 19659 6103
rect 19659 6069 19668 6103
rect 19616 6060 19668 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 10214 5958 10266 6010
rect 10278 5958 10330 6010
rect 10342 5958 10394 6010
rect 10406 5958 10458 6010
rect 10470 5958 10522 6010
rect 16214 5958 16266 6010
rect 16278 5958 16330 6010
rect 16342 5958 16394 6010
rect 16406 5958 16458 6010
rect 16470 5958 16522 6010
rect 2136 5856 2188 5908
rect 2872 5856 2924 5908
rect 3148 5856 3200 5908
rect 2596 5720 2648 5772
rect 6276 5856 6328 5908
rect 8024 5856 8076 5908
rect 11060 5856 11112 5908
rect 12440 5899 12492 5908
rect 12440 5865 12449 5899
rect 12449 5865 12483 5899
rect 12483 5865 12492 5899
rect 12440 5856 12492 5865
rect 12624 5856 12676 5908
rect 16580 5899 16632 5908
rect 16580 5865 16589 5899
rect 16589 5865 16623 5899
rect 16623 5865 16632 5899
rect 16580 5856 16632 5865
rect 16672 5856 16724 5908
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 6828 5720 6880 5772
rect 12808 5788 12860 5840
rect 2872 5516 2924 5568
rect 4804 5516 4856 5568
rect 5080 5516 5132 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 6460 5627 6512 5636
rect 6460 5593 6469 5627
rect 6469 5593 6503 5627
rect 6503 5593 6512 5627
rect 6460 5584 6512 5593
rect 6920 5584 6972 5636
rect 9036 5652 9088 5704
rect 9496 5652 9548 5704
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 10692 5652 10744 5704
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12624 5695 12676 5704
rect 12624 5661 12633 5695
rect 12633 5661 12667 5695
rect 12667 5661 12676 5695
rect 12624 5652 12676 5661
rect 18144 5763 18196 5772
rect 18144 5729 18153 5763
rect 18153 5729 18187 5763
rect 18187 5729 18196 5763
rect 18144 5720 18196 5729
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 13084 5652 13136 5704
rect 17684 5584 17736 5636
rect 8484 5516 8536 5568
rect 8576 5559 8628 5568
rect 8576 5525 8585 5559
rect 8585 5525 8619 5559
rect 8619 5525 8628 5559
rect 8576 5516 8628 5525
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 12532 5516 12584 5568
rect 12624 5516 12676 5568
rect 13728 5516 13780 5568
rect 7214 5414 7266 5466
rect 7278 5414 7330 5466
rect 7342 5414 7394 5466
rect 7406 5414 7458 5466
rect 7470 5414 7522 5466
rect 13214 5414 13266 5466
rect 13278 5414 13330 5466
rect 13342 5414 13394 5466
rect 13406 5414 13458 5466
rect 13470 5414 13522 5466
rect 19214 5414 19266 5466
rect 19278 5414 19330 5466
rect 19342 5414 19394 5466
rect 19406 5414 19458 5466
rect 19470 5414 19522 5466
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 2872 5083 2924 5092
rect 2872 5049 2881 5083
rect 2881 5049 2915 5083
rect 2915 5049 2924 5083
rect 5540 5312 5592 5364
rect 6276 5244 6328 5296
rect 7932 5312 7984 5364
rect 10048 5312 10100 5364
rect 7104 5244 7156 5296
rect 8484 5244 8536 5296
rect 3884 5176 3936 5228
rect 3976 5219 4028 5228
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 8576 5176 8628 5228
rect 2872 5040 2924 5049
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 3516 4972 3568 4981
rect 6368 5151 6420 5160
rect 6368 5117 6377 5151
rect 6377 5117 6411 5151
rect 6411 5117 6420 5151
rect 6368 5108 6420 5117
rect 8208 5040 8260 5092
rect 4804 4972 4856 5024
rect 6460 4972 6512 5024
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 9496 5244 9548 5296
rect 9956 5244 10008 5296
rect 11704 5312 11756 5364
rect 13084 5312 13136 5364
rect 9404 5176 9456 5228
rect 9680 5219 9732 5228
rect 9680 5185 9689 5219
rect 9689 5185 9723 5219
rect 9723 5185 9732 5219
rect 9680 5176 9732 5185
rect 12532 5244 12584 5296
rect 12164 5176 12216 5228
rect 12624 5176 12676 5228
rect 14464 5244 14516 5296
rect 18144 5312 18196 5364
rect 19708 5312 19760 5364
rect 19616 5244 19668 5296
rect 12624 5083 12676 5092
rect 12624 5049 12633 5083
rect 12633 5049 12667 5083
rect 12667 5049 12676 5083
rect 12624 5040 12676 5049
rect 9128 4972 9180 5024
rect 9496 4972 9548 5024
rect 13176 5151 13228 5160
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 14740 5151 14792 5160
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 20812 5176 20864 5228
rect 13360 4972 13412 5024
rect 13728 4972 13780 5024
rect 20260 5015 20312 5024
rect 20260 4981 20269 5015
rect 20269 4981 20303 5015
rect 20303 4981 20312 5015
rect 20260 4972 20312 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 10214 4870 10266 4922
rect 10278 4870 10330 4922
rect 10342 4870 10394 4922
rect 10406 4870 10458 4922
rect 10470 4870 10522 4922
rect 16214 4870 16266 4922
rect 16278 4870 16330 4922
rect 16342 4870 16394 4922
rect 16406 4870 16458 4922
rect 16470 4870 16522 4922
rect 5540 4768 5592 4820
rect 6368 4768 6420 4820
rect 9496 4811 9548 4820
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 13176 4768 13228 4820
rect 14740 4768 14792 4820
rect 14464 4700 14516 4752
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 6000 4564 6052 4616
rect 6460 4632 6512 4684
rect 8208 4564 8260 4616
rect 9036 4564 9088 4616
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9404 4564 9456 4616
rect 12992 4564 13044 4616
rect 13084 4607 13136 4616
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 3884 4496 3936 4548
rect 3976 4496 4028 4548
rect 9128 4539 9180 4548
rect 9128 4505 9137 4539
rect 9137 4505 9171 4539
rect 9171 4505 9180 4539
rect 9128 4496 9180 4505
rect 9680 4496 9732 4548
rect 20260 4564 20312 4616
rect 14188 4539 14240 4548
rect 14188 4505 14197 4539
rect 14197 4505 14231 4539
rect 14231 4505 14240 4539
rect 14188 4496 14240 4505
rect 9956 4428 10008 4480
rect 7214 4326 7266 4378
rect 7278 4326 7330 4378
rect 7342 4326 7394 4378
rect 7406 4326 7458 4378
rect 7470 4326 7522 4378
rect 13214 4326 13266 4378
rect 13278 4326 13330 4378
rect 13342 4326 13394 4378
rect 13406 4326 13458 4378
rect 13470 4326 13522 4378
rect 19214 4326 19266 4378
rect 19278 4326 19330 4378
rect 19342 4326 19394 4378
rect 19406 4326 19458 4378
rect 19470 4326 19522 4378
rect 8208 4224 8260 4276
rect 20 4088 72 4140
rect 1492 4088 1544 4140
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 9312 4088 9364 4140
rect 12164 4224 12216 4276
rect 7932 4063 7984 4072
rect 7932 4029 7941 4063
rect 7941 4029 7975 4063
rect 7975 4029 7984 4063
rect 7932 4020 7984 4029
rect 8208 4063 8260 4072
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 8208 4020 8260 4029
rect 8668 4020 8720 4072
rect 9404 4020 9456 4072
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 7656 3884 7708 3893
rect 9220 3884 9272 3936
rect 9956 3884 10008 3936
rect 12624 4156 12676 4208
rect 11980 4063 12032 4072
rect 11980 4029 11989 4063
rect 11989 4029 12023 4063
rect 12023 4029 12032 4063
rect 11980 4020 12032 4029
rect 10692 3952 10744 4004
rect 13084 4088 13136 4140
rect 20628 4020 20680 4072
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 11888 3884 11940 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 12716 3884 12768 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 10214 3782 10266 3834
rect 10278 3782 10330 3834
rect 10342 3782 10394 3834
rect 10406 3782 10458 3834
rect 10470 3782 10522 3834
rect 16214 3782 16266 3834
rect 16278 3782 16330 3834
rect 16342 3782 16394 3834
rect 16406 3782 16458 3834
rect 16470 3782 16522 3834
rect 6000 3723 6052 3732
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 7656 3680 7708 3732
rect 8208 3680 8260 3732
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 6920 3519 6972 3528
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 8300 3476 8352 3528
rect 3884 3408 3936 3460
rect 4528 3451 4580 3460
rect 4528 3417 4537 3451
rect 4537 3417 4571 3451
rect 4571 3417 4580 3451
rect 4528 3408 4580 3417
rect 5080 3408 5132 3460
rect 8116 3340 8168 3392
rect 9404 3476 9456 3528
rect 10600 3680 10652 3732
rect 11888 3680 11940 3732
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 11980 3519 12032 3528
rect 9128 3451 9180 3460
rect 9128 3417 9137 3451
rect 9137 3417 9171 3451
rect 9171 3417 9180 3451
rect 9128 3408 9180 3417
rect 9220 3451 9272 3460
rect 9220 3417 9229 3451
rect 9229 3417 9263 3451
rect 9263 3417 9272 3451
rect 9220 3408 9272 3417
rect 9312 3340 9364 3392
rect 9956 3340 10008 3392
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 12532 3476 12584 3528
rect 11796 3340 11848 3392
rect 11888 3383 11940 3392
rect 11888 3349 11897 3383
rect 11897 3349 11931 3383
rect 11931 3349 11940 3383
rect 11888 3340 11940 3349
rect 12348 3340 12400 3392
rect 12532 3340 12584 3392
rect 7214 3238 7266 3290
rect 7278 3238 7330 3290
rect 7342 3238 7394 3290
rect 7406 3238 7458 3290
rect 7470 3238 7522 3290
rect 13214 3238 13266 3290
rect 13278 3238 13330 3290
rect 13342 3238 13394 3290
rect 13406 3238 13458 3290
rect 13470 3238 13522 3290
rect 19214 3238 19266 3290
rect 19278 3238 19330 3290
rect 19342 3238 19394 3290
rect 19406 3238 19458 3290
rect 19470 3238 19522 3290
rect 4528 3136 4580 3188
rect 6920 3136 6972 3188
rect 7932 3136 7984 3188
rect 10416 3136 10468 3188
rect 10692 3136 10744 3188
rect 3516 3068 3568 3120
rect 5080 3068 5132 3120
rect 8668 3000 8720 3052
rect 9312 3000 9364 3052
rect 3884 2932 3936 2984
rect 9680 2932 9732 2984
rect 11796 3136 11848 3188
rect 11980 3136 12032 3188
rect 12072 3136 12124 3188
rect 11796 3043 11848 3052
rect 11796 3009 11800 3043
rect 11800 3009 11834 3043
rect 11834 3009 11848 3043
rect 11796 3000 11848 3009
rect 12532 3068 12584 3120
rect 14556 3136 14608 3188
rect 14924 3068 14976 3120
rect 11612 2907 11664 2916
rect 11612 2873 11621 2907
rect 11621 2873 11655 2907
rect 11655 2873 11664 2907
rect 11612 2864 11664 2873
rect 12624 2975 12676 2984
rect 12624 2941 12633 2975
rect 12633 2941 12667 2975
rect 12667 2941 12676 2975
rect 12624 2932 12676 2941
rect 14188 2975 14240 2984
rect 14188 2941 14197 2975
rect 14197 2941 14231 2975
rect 14231 2941 14240 2975
rect 14188 2932 14240 2941
rect 12716 2796 12768 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 10214 2694 10266 2746
rect 10278 2694 10330 2746
rect 10342 2694 10394 2746
rect 10406 2694 10458 2746
rect 10470 2694 10522 2746
rect 16214 2694 16266 2746
rect 16278 2694 16330 2746
rect 16342 2694 16394 2746
rect 16406 2694 16458 2746
rect 16470 2694 16522 2746
rect 8760 2592 8812 2644
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 14188 2592 14240 2644
rect 9680 2456 9732 2508
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 12532 2388 12584 2440
rect 15200 2388 15252 2440
rect 15568 2363 15620 2372
rect 15568 2329 15577 2363
rect 15577 2329 15611 2363
rect 15611 2329 15620 2363
rect 15568 2320 15620 2329
rect 7214 2150 7266 2202
rect 7278 2150 7330 2202
rect 7342 2150 7394 2202
rect 7406 2150 7458 2202
rect 7470 2150 7522 2202
rect 13214 2150 13266 2202
rect 13278 2150 13330 2202
rect 13342 2150 13394 2202
rect 13406 2150 13458 2202
rect 13470 2150 13522 2202
rect 19214 2150 19266 2202
rect 19278 2150 19330 2202
rect 19342 2150 19394 2202
rect 19406 2150 19458 2202
rect 19470 2150 19522 2202
<< metal2 >>
rect 3238 23262 3294 24062
rect 8390 23262 8446 24062
rect 13542 23262 13598 24062
rect 18694 23262 18750 24062
rect 3252 22094 3280 23262
rect 3252 22066 3372 22094
rect 3146 21856 3202 21865
rect 3146 21791 3202 21800
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 2136 17740 2188 17746
rect 2136 17682 2188 17688
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1596 16522 1624 17614
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 1584 16516 1636 16522
rect 1584 16458 1636 16464
rect 952 16425 980 16458
rect 938 16416 994 16425
rect 938 16351 994 16360
rect 1596 16182 1624 16458
rect 1584 16176 1636 16182
rect 1584 16118 1636 16124
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14618 1532 14758
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1688 14498 1716 16594
rect 1872 15416 1900 17682
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1964 16250 1992 17138
rect 2148 16590 2176 17682
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1952 15428 2004 15434
rect 1872 15388 1952 15416
rect 1952 15370 2004 15376
rect 1964 14958 1992 15370
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1688 14470 1808 14498
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 1688 12986 1716 13194
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 10985 1440 11698
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10266 1624 10406
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9586 1716 9862
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8498 1716 8774
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 6914 1624 7278
rect 1504 6886 1624 6914
rect 1780 6914 1808 14470
rect 1964 14346 1992 14894
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 2056 14074 2084 16050
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 12238 1900 13806
rect 2056 13394 2084 14010
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2148 12646 2176 14758
rect 2332 14618 2360 15030
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2792 13326 2820 14350
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2320 13184 2372 13190
rect 2884 13172 2912 18566
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2976 17134 3004 17478
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 3068 16522 3096 16934
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 3160 16266 3188 21791
rect 3344 21554 3372 22066
rect 7214 21788 7522 21797
rect 7214 21786 7220 21788
rect 7276 21786 7300 21788
rect 7356 21786 7380 21788
rect 7436 21786 7460 21788
rect 7516 21786 7522 21788
rect 7276 21734 7278 21786
rect 7458 21734 7460 21786
rect 7214 21732 7220 21734
rect 7276 21732 7300 21734
rect 7356 21732 7380 21734
rect 7436 21732 7460 21734
rect 7516 21732 7522 21734
rect 7214 21723 7522 21732
rect 3332 21548 3384 21554
rect 3332 21490 3384 21496
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4080 19854 4108 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4080 19514 4108 19654
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 3252 18970 3280 19110
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 4080 18952 4108 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18970 4660 19314
rect 4160 18964 4212 18970
rect 4080 18924 4160 18952
rect 4080 17542 4108 18924
rect 4160 18906 4212 18912
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4724 17746 4752 18158
rect 4816 17746 4844 21286
rect 8404 20942 8432 23262
rect 13556 22094 13584 23262
rect 13556 22066 13860 22094
rect 13214 21788 13522 21797
rect 13214 21786 13220 21788
rect 13276 21786 13300 21788
rect 13356 21786 13380 21788
rect 13436 21786 13460 21788
rect 13516 21786 13522 21788
rect 13276 21734 13278 21786
rect 13458 21734 13460 21786
rect 13214 21732 13220 21734
rect 13276 21732 13300 21734
rect 13356 21732 13380 21734
rect 13436 21732 13460 21734
rect 13516 21732 13522 21734
rect 13214 21723 13522 21732
rect 13832 21554 13860 22066
rect 18708 21554 18736 23262
rect 19214 21788 19522 21797
rect 19214 21786 19220 21788
rect 19276 21786 19300 21788
rect 19356 21786 19380 21788
rect 19436 21786 19460 21788
rect 19516 21786 19522 21788
rect 19276 21734 19278 21786
rect 19458 21734 19460 21786
rect 19214 21732 19220 21734
rect 19276 21732 19300 21734
rect 19356 21732 19380 21734
rect 19436 21732 19460 21734
rect 19516 21732 19522 21734
rect 19214 21723 19522 21732
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 10214 21244 10522 21253
rect 10214 21242 10220 21244
rect 10276 21242 10300 21244
rect 10356 21242 10380 21244
rect 10436 21242 10460 21244
rect 10516 21242 10522 21244
rect 10276 21190 10278 21242
rect 10458 21190 10460 21242
rect 10214 21188 10220 21190
rect 10276 21188 10300 21190
rect 10356 21188 10380 21190
rect 10436 21188 10460 21190
rect 10516 21188 10522 21190
rect 10214 21179 10522 21188
rect 12452 21146 12480 21286
rect 14384 21146 14412 21422
rect 16214 21244 16522 21253
rect 16214 21242 16220 21244
rect 16276 21242 16300 21244
rect 16356 21242 16380 21244
rect 16436 21242 16460 21244
rect 16516 21242 16522 21244
rect 16276 21190 16278 21242
rect 16458 21190 16460 21242
rect 16214 21188 16220 21190
rect 16276 21188 16300 21190
rect 16356 21188 16380 21190
rect 16436 21188 16460 21190
rect 16516 21188 16522 21190
rect 16214 21179 16522 21188
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4908 20466 4936 20742
rect 7024 20466 7052 20878
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4816 17610 4844 17682
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 5184 17338 5212 18770
rect 5736 18766 5764 19110
rect 5828 18902 5856 20198
rect 6012 19854 6040 20402
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6564 19854 6592 20198
rect 7116 20058 7144 20878
rect 8760 20868 8812 20874
rect 8760 20810 8812 20816
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 8300 20800 8352 20806
rect 8300 20742 8352 20748
rect 7214 20700 7522 20709
rect 7214 20698 7220 20700
rect 7276 20698 7300 20700
rect 7356 20698 7380 20700
rect 7436 20698 7460 20700
rect 7516 20698 7522 20700
rect 7276 20646 7278 20698
rect 7458 20646 7460 20698
rect 7214 20644 7220 20646
rect 7276 20644 7300 20646
rect 7356 20644 7380 20646
rect 7436 20644 7460 20646
rect 7516 20644 7522 20646
rect 7214 20635 7522 20644
rect 7576 20534 7604 20742
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 8312 20398 8340 20742
rect 8772 20602 8800 20810
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 10336 20466 10364 20742
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6460 19848 6512 19854
rect 6460 19790 6512 19796
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6288 19514 6316 19790
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6380 19514 6408 19654
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5920 18834 5948 19314
rect 6288 18970 6316 19314
rect 6472 18970 6500 19790
rect 7214 19612 7522 19621
rect 7214 19610 7220 19612
rect 7276 19610 7300 19612
rect 7356 19610 7380 19612
rect 7436 19610 7460 19612
rect 7516 19610 7522 19612
rect 7276 19558 7278 19610
rect 7458 19558 7460 19610
rect 7214 19556 7220 19558
rect 7276 19556 7300 19558
rect 7356 19556 7380 19558
rect 7436 19556 7460 19558
rect 7516 19556 7522 19558
rect 7214 19547 7522 19556
rect 8312 19378 8340 20334
rect 10152 20058 10180 20402
rect 10214 20156 10522 20165
rect 10214 20154 10220 20156
rect 10276 20154 10300 20156
rect 10356 20154 10380 20156
rect 10436 20154 10460 20156
rect 10516 20154 10522 20156
rect 10276 20102 10278 20154
rect 10458 20102 10460 20154
rect 10214 20100 10220 20102
rect 10276 20100 10300 20102
rect 10356 20100 10380 20102
rect 10436 20100 10460 20102
rect 10516 20100 10522 20102
rect 10214 20091 10522 20100
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 10796 19854 10824 20742
rect 11624 20602 11652 20810
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 12544 20534 12572 20742
rect 10876 20528 10928 20534
rect 10876 20470 10928 20476
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 7852 18902 7880 19110
rect 8588 18970 8616 19246
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5920 18698 5948 18770
rect 5908 18692 5960 18698
rect 5908 18634 5960 18640
rect 7214 18524 7522 18533
rect 7214 18522 7220 18524
rect 7276 18522 7300 18524
rect 7356 18522 7380 18524
rect 7436 18522 7460 18524
rect 7516 18522 7522 18524
rect 7276 18470 7278 18522
rect 7458 18470 7460 18522
rect 7214 18468 7220 18470
rect 7276 18468 7300 18470
rect 7356 18468 7380 18470
rect 7436 18468 7460 18470
rect 7516 18468 7522 18470
rect 7214 18459 7522 18468
rect 7852 18408 7880 18838
rect 9324 18834 9352 19450
rect 10796 19378 10824 19790
rect 10888 19378 10916 20470
rect 12452 19854 12480 20470
rect 12636 20262 12664 20878
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 13214 20700 13522 20709
rect 13214 20698 13220 20700
rect 13276 20698 13300 20700
rect 13356 20698 13380 20700
rect 13436 20698 13460 20700
rect 13516 20698 13522 20700
rect 13276 20646 13278 20698
rect 13458 20646 13460 20698
rect 13214 20644 13220 20646
rect 13276 20644 13300 20646
rect 13356 20644 13380 20646
rect 13436 20644 13460 20646
rect 13516 20644 13522 20646
rect 13214 20635 13522 20644
rect 14200 20534 14228 20742
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12636 20058 12664 20198
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9324 18426 9352 18770
rect 9312 18420 9364 18426
rect 7852 18380 8064 18408
rect 8036 18290 8064 18380
rect 9312 18362 9364 18368
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 9324 17882 9352 18362
rect 10060 18290 10088 19314
rect 11164 19174 11192 19654
rect 11808 19242 11836 19722
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 19446 12296 19654
rect 12912 19446 12940 19994
rect 13740 19854 13768 20402
rect 14200 19854 14228 20470
rect 15212 20262 15240 20810
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13214 19612 13522 19621
rect 13214 19610 13220 19612
rect 13276 19610 13300 19612
rect 13356 19610 13380 19612
rect 13436 19610 13460 19612
rect 13516 19610 13522 19612
rect 13276 19558 13278 19610
rect 13458 19558 13460 19610
rect 13214 19556 13220 19558
rect 13276 19556 13300 19558
rect 13356 19556 13380 19558
rect 13436 19556 13460 19558
rect 13516 19556 13522 19558
rect 13214 19547 13522 19556
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12900 19440 12952 19446
rect 12900 19382 12952 19388
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 10214 19068 10522 19077
rect 10214 19066 10220 19068
rect 10276 19066 10300 19068
rect 10356 19066 10380 19068
rect 10436 19066 10460 19068
rect 10516 19066 10522 19068
rect 10276 19014 10278 19066
rect 10458 19014 10460 19066
rect 10214 19012 10220 19014
rect 10276 19012 10300 19014
rect 10356 19012 10380 19014
rect 10436 19012 10460 19014
rect 10516 19012 10522 19014
rect 10214 19003 10522 19012
rect 10796 18970 10824 19110
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 11808 18698 11836 19178
rect 12912 18970 12940 19382
rect 13832 19174 13860 19722
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19514 14136 19654
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 11796 18692 11848 18698
rect 11796 18634 11848 18640
rect 12452 18426 12480 18906
rect 13214 18524 13522 18533
rect 13214 18522 13220 18524
rect 13276 18522 13300 18524
rect 13356 18522 13380 18524
rect 13436 18522 13460 18524
rect 13516 18522 13522 18524
rect 13276 18470 13278 18522
rect 13458 18470 13460 18522
rect 13214 18468 13220 18470
rect 13276 18468 13300 18470
rect 13356 18468 13380 18470
rect 13436 18468 13460 18470
rect 13516 18468 13522 18470
rect 13214 18459 13522 18468
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9324 17678 9352 17818
rect 9784 17762 9812 18022
rect 9416 17734 9812 17762
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 5828 17542 5856 17614
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 3608 17264 3660 17270
rect 3608 17206 3660 17212
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3528 16794 3556 16934
rect 3620 16794 3648 17206
rect 5184 17202 5212 17274
rect 5828 17202 5856 17478
rect 6564 17338 6592 17546
rect 9416 17542 9444 17734
rect 9784 17610 9812 17734
rect 9772 17604 9824 17610
rect 9772 17546 9824 17552
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 7214 17436 7522 17445
rect 7214 17434 7220 17436
rect 7276 17434 7300 17436
rect 7356 17434 7380 17436
rect 7436 17434 7460 17436
rect 7516 17434 7522 17436
rect 7276 17382 7278 17434
rect 7458 17382 7460 17434
rect 7214 17380 7220 17382
rect 7276 17380 7300 17382
rect 7356 17380 7380 17382
rect 7436 17380 7460 17382
rect 7516 17380 7522 17382
rect 7214 17371 7522 17380
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 4620 16992 4672 16998
rect 3712 16918 4016 16946
rect 4620 16934 4672 16940
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3160 16238 3280 16266
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2320 13126 2372 13132
rect 2792 13144 2912 13172
rect 2332 12986 2360 13126
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 2148 12170 2176 12582
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 2148 11898 2176 12106
rect 2516 11898 2544 12718
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2332 10810 2360 10950
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2516 10742 2544 11834
rect 2792 11218 2820 13144
rect 2976 12918 3004 13194
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12442 2912 12718
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 3160 12306 3188 13398
rect 3252 12434 3280 16238
rect 3344 15570 3372 16390
rect 3528 15910 3556 16730
rect 3712 16658 3740 16918
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3896 16590 3924 16730
rect 3988 16658 4016 16918
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3896 16454 3924 16526
rect 4632 16522 4660 16934
rect 5000 16794 5028 17138
rect 7576 17134 7604 17478
rect 8680 17338 8708 17478
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 9508 17134 9536 17478
rect 10060 17202 10088 18226
rect 10214 17980 10522 17989
rect 10214 17978 10220 17980
rect 10276 17978 10300 17980
rect 10356 17978 10380 17980
rect 10436 17978 10460 17980
rect 10516 17978 10522 17980
rect 10276 17926 10278 17978
rect 10458 17926 10460 17978
rect 10214 17924 10220 17926
rect 10276 17924 10300 17926
rect 10356 17924 10380 17926
rect 10436 17924 10460 17926
rect 10516 17924 10522 17926
rect 10214 17915 10522 17924
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10336 17338 10364 17478
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10520 17202 10548 17478
rect 11072 17202 11100 17478
rect 12452 17338 12480 18362
rect 13740 17882 13768 18906
rect 14568 18902 14596 19382
rect 15028 19378 15056 20198
rect 15212 20058 15240 20198
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 14108 18086 14136 18634
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14200 18290 14228 18566
rect 14384 18426 14412 18566
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13214 17436 13522 17445
rect 13214 17434 13220 17436
rect 13276 17434 13300 17436
rect 13356 17434 13380 17436
rect 13436 17434 13460 17436
rect 13516 17434 13522 17436
rect 13276 17382 13278 17434
rect 13458 17382 13460 17434
rect 13214 17380 13220 17382
rect 13276 17380 13300 17382
rect 13356 17380 13380 17382
rect 13436 17380 13460 17382
rect 13516 17380 13522 17382
rect 13214 17371 13522 17380
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10508 17196 10560 17202
rect 11060 17196 11112 17202
rect 10560 17156 10640 17184
rect 10508 17138 10560 17144
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5552 16590 5580 16934
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 7116 16454 7144 16934
rect 8588 16658 8616 17070
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12918 3372 13262
rect 3528 13258 3556 15846
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14618 3740 14894
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3804 14482 3832 15302
rect 3896 14958 3924 15438
rect 3988 15434 4016 16390
rect 7214 16348 7522 16357
rect 7214 16346 7220 16348
rect 7276 16346 7300 16348
rect 7356 16346 7380 16348
rect 7436 16346 7460 16348
rect 7516 16346 7522 16348
rect 7276 16294 7278 16346
rect 7458 16294 7460 16346
rect 7214 16292 7220 16294
rect 7276 16292 7300 16294
rect 7356 16292 7380 16294
rect 7436 16292 7460 16294
rect 7516 16292 7522 16294
rect 7214 16283 7522 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 4172 15094 4200 15438
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 14482 4752 15302
rect 4908 15162 4936 15438
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 5276 14618 5304 15030
rect 6196 14958 6224 15370
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 5920 14618 5948 14894
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 6288 13530 6316 14418
rect 6380 14414 6408 15506
rect 6644 15428 6696 15434
rect 6644 15370 6696 15376
rect 6656 15162 6684 15370
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7214 15260 7522 15269
rect 7214 15258 7220 15260
rect 7276 15258 7300 15260
rect 7356 15258 7380 15260
rect 7436 15258 7460 15260
rect 7516 15258 7522 15260
rect 7276 15206 7278 15258
rect 7458 15206 7460 15258
rect 7214 15204 7220 15206
rect 7276 15204 7300 15206
rect 7356 15204 7380 15206
rect 7436 15204 7460 15206
rect 7516 15204 7522 15206
rect 7214 15195 7522 15204
rect 7668 15162 7696 15302
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 6472 14618 6500 14962
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6748 14618 6776 14894
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14618 7788 14758
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6380 14006 6408 14350
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 7024 13938 7052 14214
rect 7214 14172 7522 14181
rect 7214 14170 7220 14172
rect 7276 14170 7300 14172
rect 7356 14170 7380 14172
rect 7436 14170 7460 14172
rect 7516 14170 7522 14172
rect 7276 14118 7278 14170
rect 7458 14118 7460 14170
rect 7214 14116 7220 14118
rect 7276 14116 7300 14118
rect 7356 14116 7380 14118
rect 7436 14116 7460 14118
rect 7516 14116 7522 14118
rect 7214 14107 7522 14116
rect 7760 14074 7788 14554
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7852 14006 7880 16390
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 8036 15026 8064 15370
rect 8588 15026 8616 16594
rect 8024 15020 8076 15026
rect 8024 14962 8076 14968
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8496 14074 8524 14962
rect 8588 14618 8616 14962
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 7840 14000 7892 14006
rect 7760 13948 7840 13954
rect 7760 13942 7892 13948
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7760 13926 7880 13942
rect 8392 13932 8444 13938
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 3332 12912 3384 12918
rect 3384 12860 3924 12866
rect 3332 12854 3924 12860
rect 3344 12838 3924 12854
rect 3252 12406 3372 12434
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3252 11286 3280 12174
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2516 10130 2544 10678
rect 2700 10266 2728 10950
rect 2884 10266 2912 11086
rect 3252 10742 3280 11222
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2516 9722 2544 10066
rect 3252 10062 3280 10678
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2240 9178 2268 9318
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2228 7948 2280 7954
rect 2228 7890 2280 7896
rect 1780 6886 2176 6914
rect 1504 6730 1532 6886
rect 1492 6724 1544 6730
rect 1492 6666 1544 6672
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1504 4146 1532 6666
rect 2148 5914 2176 6886
rect 2240 6866 2268 7890
rect 2424 7478 2452 8230
rect 2516 7954 2544 9658
rect 3344 9178 3372 12406
rect 3896 12374 3924 12838
rect 4264 12696 4292 13194
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4540 12986 4568 13126
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 5736 12918 5764 13194
rect 6656 12986 6684 13262
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 4436 12776 4488 12782
rect 4488 12736 4752 12764
rect 4436 12718 4488 12724
rect 4080 12668 4292 12696
rect 4080 12442 4108 12668
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4724 12442 4752 12736
rect 5736 12714 5764 12854
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4540 11898 4568 12174
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5460 11218 5488 12038
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 3988 10810 4016 11018
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3988 10266 4016 10746
rect 4540 10674 4568 10950
rect 4632 10690 4660 11018
rect 4724 10810 4752 11018
rect 5356 11008 5408 11014
rect 5460 10996 5488 11154
rect 5724 11008 5776 11014
rect 5460 10968 5580 10996
rect 5356 10950 5408 10956
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4528 10668 4580 10674
rect 4632 10662 4752 10690
rect 4528 10610 4580 10616
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4080 9926 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10130 4660 10474
rect 4724 10470 4752 10662
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4724 9994 4752 10406
rect 4816 10266 4844 10542
rect 5276 10266 5304 10746
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3804 8634 3832 9590
rect 4816 9382 4844 10066
rect 5276 9994 5304 10202
rect 5368 10130 5396 10950
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 10266 5488 10406
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5092 9450 5120 9862
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 8634 4384 8774
rect 4448 8634 4476 8978
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4724 8498 4752 8910
rect 4816 8634 4844 9318
rect 5092 9042 5120 9386
rect 5276 9042 5304 9930
rect 5552 9654 5580 10968
rect 5724 10950 5776 10956
rect 5736 10742 5764 10950
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5736 10266 5764 10678
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 6368 10192 6420 10198
rect 6368 10134 6420 10140
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 5000 8566 5028 8774
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4160 8424 4212 8430
rect 3988 8384 4160 8412
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 8090 3924 8230
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3160 7750 3188 7890
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3712 7546 3740 7754
rect 3988 7750 4016 8384
rect 4160 8366 4212 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4816 7818 4844 7890
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 4080 7546 4108 7754
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2608 5778 2636 6054
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2792 5370 2820 6258
rect 2884 5914 2912 6258
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5914 3188 6054
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2884 5098 2912 5510
rect 3988 5234 4016 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4816 5574 4844 7754
rect 5092 7410 5120 8978
rect 5276 8634 5304 8978
rect 5736 8634 5764 10066
rect 6092 9988 6144 9994
rect 6092 9930 6144 9936
rect 6104 9586 6132 9930
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5184 7410 5212 8230
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5368 7410 5396 8026
rect 5552 7954 5580 8230
rect 5828 8090 5856 8230
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5552 7410 5580 7890
rect 5920 7818 5948 8366
rect 6104 7886 6132 9522
rect 6288 9178 6316 9590
rect 6380 9586 6408 10134
rect 6472 9994 6500 12650
rect 6748 12434 6776 13670
rect 6932 13394 6960 13874
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6932 12850 6960 13330
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7024 12714 7052 13194
rect 7214 13084 7522 13093
rect 7214 13082 7220 13084
rect 7276 13082 7300 13084
rect 7356 13082 7380 13084
rect 7436 13082 7460 13084
rect 7516 13082 7522 13084
rect 7276 13030 7278 13082
rect 7458 13030 7460 13082
rect 7214 13028 7220 13030
rect 7276 13028 7300 13030
rect 7356 13028 7380 13030
rect 7436 13028 7460 13030
rect 7516 13028 7522 13030
rect 7214 13019 7522 13028
rect 7760 12850 7788 13926
rect 8392 13874 8444 13880
rect 8404 13530 8432 13874
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8496 12918 8524 14010
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8588 13190 8616 13874
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 8404 12434 8432 12718
rect 8484 12436 8536 12442
rect 6748 12406 6868 12434
rect 8404 12406 8484 12434
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6564 9722 6592 10610
rect 6656 10198 6684 10610
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6748 9586 6776 10406
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6196 8634 6224 9114
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6288 8498 6316 9114
rect 6380 8974 6408 9522
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6196 8022 6224 8434
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 6012 7546 6040 7822
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 6104 7342 6132 7822
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7546 6224 7686
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6288 7410 6316 8434
rect 6656 7818 6684 9318
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6748 8090 6776 8842
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6748 7954 6776 8026
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6288 7002 6316 7346
rect 6656 7206 6684 7754
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6288 6458 6316 6938
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6288 5914 6316 6394
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6840 5778 6868 12406
rect 8484 12378 8536 12384
rect 7214 11996 7522 12005
rect 7214 11994 7220 11996
rect 7276 11994 7300 11996
rect 7356 11994 7380 11996
rect 7436 11994 7460 11996
rect 7516 11994 7522 11996
rect 7276 11942 7278 11994
rect 7458 11942 7460 11994
rect 7214 11940 7220 11942
rect 7276 11940 7300 11942
rect 7356 11940 7380 11942
rect 7436 11940 7460 11942
rect 7516 11940 7522 11942
rect 7214 11931 7522 11940
rect 8588 11234 8616 13126
rect 8404 11206 8616 11234
rect 8404 11082 8432 11206
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 7214 10908 7522 10917
rect 7214 10906 7220 10908
rect 7276 10906 7300 10908
rect 7356 10906 7380 10908
rect 7436 10906 7460 10908
rect 7516 10906 7522 10908
rect 7276 10854 7278 10906
rect 7458 10854 7460 10906
rect 7214 10852 7220 10854
rect 7276 10852 7300 10854
rect 7356 10852 7380 10854
rect 7436 10852 7460 10854
rect 7516 10852 7522 10854
rect 7214 10843 7522 10852
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6932 9586 6960 10542
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 10130 7420 10406
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 7760 9994 7788 10610
rect 8312 10606 8340 10950
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7214 9820 7522 9829
rect 7214 9818 7220 9820
rect 7276 9818 7300 9820
rect 7356 9818 7380 9820
rect 7436 9818 7460 9820
rect 7516 9818 7522 9820
rect 7276 9766 7278 9818
rect 7458 9766 7460 9818
rect 7214 9764 7220 9766
rect 7276 9764 7300 9766
rect 7356 9764 7380 9766
rect 7436 9764 7460 9766
rect 7516 9764 7522 9766
rect 7214 9755 7522 9764
rect 7760 9722 7788 9930
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 8220 9654 8248 9998
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 6932 9110 6960 9522
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7760 9042 7788 9522
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7944 8974 7972 9522
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7024 7886 7052 8774
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7546 6960 7754
rect 7012 7744 7064 7750
rect 7116 7698 7144 8774
rect 7214 8732 7522 8741
rect 7214 8730 7220 8732
rect 7276 8730 7300 8732
rect 7356 8730 7380 8732
rect 7436 8730 7460 8732
rect 7516 8730 7522 8732
rect 7276 8678 7278 8730
rect 7458 8678 7460 8730
rect 7214 8676 7220 8678
rect 7276 8676 7300 8678
rect 7356 8676 7380 8678
rect 7436 8676 7460 8678
rect 7516 8676 7522 8678
rect 7214 8667 7522 8676
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7886 7236 8230
rect 7300 8090 7328 8366
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7484 7834 7512 8502
rect 7576 8090 7604 8910
rect 8128 8838 8156 9522
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7668 8090 7696 8774
rect 7760 8362 7788 8774
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 8090 7880 8230
rect 8220 8090 8248 9590
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8312 9178 8340 9454
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8404 8412 8432 11018
rect 8496 10266 8524 11086
rect 8680 11082 8708 16934
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 10060 15314 10088 17138
rect 10214 16892 10522 16901
rect 10214 16890 10220 16892
rect 10276 16890 10300 16892
rect 10356 16890 10380 16892
rect 10436 16890 10460 16892
rect 10516 16890 10522 16892
rect 10276 16838 10278 16890
rect 10458 16838 10460 16890
rect 10214 16836 10220 16838
rect 10276 16836 10300 16838
rect 10356 16836 10380 16838
rect 10436 16836 10460 16838
rect 10516 16836 10522 16838
rect 10214 16827 10522 16836
rect 10612 16182 10640 17156
rect 11060 17138 11112 17144
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10888 16794 10916 16934
rect 12360 16794 12388 17138
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10980 16538 11008 16594
rect 10980 16510 11100 16538
rect 10600 16176 10652 16182
rect 10652 16136 10732 16164
rect 10600 16118 10652 16124
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10152 15416 10180 16050
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10214 15804 10522 15813
rect 10214 15802 10220 15804
rect 10276 15802 10300 15804
rect 10356 15802 10380 15804
rect 10436 15802 10460 15804
rect 10516 15802 10522 15804
rect 10276 15750 10278 15802
rect 10458 15750 10460 15802
rect 10214 15748 10220 15750
rect 10276 15748 10300 15750
rect 10356 15748 10380 15750
rect 10436 15748 10460 15750
rect 10516 15748 10522 15750
rect 10214 15739 10522 15748
rect 10612 15706 10640 15846
rect 10704 15706 10732 16136
rect 11072 15910 11100 16510
rect 12452 16250 12480 17274
rect 13740 17270 13768 17818
rect 14108 17270 14136 18022
rect 14200 17882 14228 18226
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14384 17678 14412 18362
rect 14476 18358 14504 18566
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14660 18086 14688 18362
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 14096 17264 14148 17270
rect 14096 17206 14148 17212
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12820 16182 12848 16934
rect 13740 16794 13768 17206
rect 15212 16794 15240 19178
rect 15396 18834 15424 19654
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15396 18222 15424 18770
rect 15488 18766 15516 20878
rect 15580 20262 15608 20878
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15580 19854 15608 20198
rect 16214 20156 16522 20165
rect 16214 20154 16220 20156
rect 16276 20154 16300 20156
rect 16356 20154 16380 20156
rect 16436 20154 16460 20156
rect 16516 20154 16522 20156
rect 16276 20102 16278 20154
rect 16458 20102 16460 20154
rect 16214 20100 16220 20102
rect 16276 20100 16300 20102
rect 16356 20100 16380 20102
rect 16436 20100 16460 20102
rect 16516 20100 16522 20102
rect 16214 20091 16522 20100
rect 16960 20058 16988 20470
rect 17328 20466 17356 20878
rect 17788 20534 17816 21490
rect 17960 21480 18012 21486
rect 17960 21422 18012 21428
rect 17972 20874 18000 21422
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18064 21146 18092 21286
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17328 20058 17356 20402
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 16120 19780 16172 19786
rect 16120 19722 16172 19728
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15396 17882 15424 18158
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 15396 17338 15424 17818
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10704 15434 10732 15642
rect 11072 15502 11100 15846
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10232 15428 10284 15434
rect 10152 15388 10232 15416
rect 10232 15370 10284 15376
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 9232 15162 9260 15302
rect 10060 15286 10180 15314
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 10152 15026 10180 15286
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10152 14006 10180 14962
rect 10244 14958 10272 15370
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10214 14716 10522 14725
rect 10214 14714 10220 14716
rect 10276 14714 10300 14716
rect 10356 14714 10380 14716
rect 10436 14714 10460 14716
rect 10516 14714 10522 14716
rect 10276 14662 10278 14714
rect 10458 14662 10460 14714
rect 10214 14660 10220 14662
rect 10276 14660 10300 14662
rect 10356 14660 10380 14662
rect 10436 14660 10460 14662
rect 10516 14660 10522 14662
rect 10214 14651 10522 14660
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8772 13394 8800 13670
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 9140 13258 9168 13874
rect 10508 13864 10560 13870
rect 10560 13812 10640 13818
rect 10508 13806 10640 13812
rect 10520 13790 10640 13806
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9508 12986 9536 13194
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 9364 8524 9454
rect 8576 9376 8628 9382
rect 8496 9336 8576 9364
rect 8496 9110 8524 9336
rect 8576 9318 8628 9324
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8484 8424 8536 8430
rect 8404 8384 8484 8412
rect 8484 8366 8536 8372
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7576 7834 7604 7890
rect 7484 7806 7604 7834
rect 7064 7692 7144 7698
rect 7012 7686 7144 7692
rect 7024 7670 7144 7686
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 7024 7206 7052 7670
rect 7214 7644 7522 7653
rect 7214 7642 7220 7644
rect 7276 7642 7300 7644
rect 7356 7642 7380 7644
rect 7436 7642 7460 7644
rect 7516 7642 7522 7644
rect 7276 7590 7278 7642
rect 7458 7590 7460 7642
rect 7214 7588 7220 7590
rect 7276 7588 7300 7590
rect 7356 7588 7380 7590
rect 7436 7588 7460 7590
rect 7516 7588 7522 7590
rect 7214 7579 7522 7588
rect 7104 7472 7156 7478
rect 7576 7460 7604 7806
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7156 7432 7604 7460
rect 7104 7414 7156 7420
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7116 7018 7144 7414
rect 6932 6990 7144 7018
rect 6932 6322 6960 6990
rect 7214 6556 7522 6565
rect 7214 6554 7220 6556
rect 7276 6554 7300 6556
rect 7356 6554 7380 6556
rect 7436 6554 7460 6556
rect 7516 6554 7522 6556
rect 7276 6502 7278 6554
rect 7458 6502 7460 6554
rect 7214 6500 7220 6502
rect 7276 6500 7300 6502
rect 7356 6500 7380 6502
rect 7436 6500 7460 6502
rect 7516 6500 7522 6502
rect 7214 6491 7522 6500
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7576 6322 7604 6394
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6932 5642 6960 6258
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 20 4140 72 4146
rect 20 4082 72 4088
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 32 800 60 4082
rect 3528 3126 3556 4966
rect 3896 4554 3924 5170
rect 3988 4554 4016 5170
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4816 4622 4844 4966
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 3884 4548 3936 4554
rect 3884 4490 3936 4496
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3896 3466 3924 4490
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5092 3466 5120 5510
rect 5552 5370 5580 5510
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5552 4826 5580 5306
rect 6276 5296 6328 5302
rect 6274 5264 6276 5273
rect 6328 5264 6330 5273
rect 6274 5199 6330 5208
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4826 6408 5102
rect 6472 5030 6500 5578
rect 7214 5468 7522 5477
rect 7214 5466 7220 5468
rect 7276 5466 7300 5468
rect 7356 5466 7380 5468
rect 7436 5466 7460 5468
rect 7516 5466 7522 5468
rect 7276 5414 7278 5466
rect 7458 5414 7460 5466
rect 7214 5412 7220 5414
rect 7276 5412 7300 5414
rect 7356 5412 7380 5414
rect 7436 5412 7460 5414
rect 7516 5412 7522 5414
rect 7214 5403 7522 5412
rect 7944 5370 7972 7754
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 5914 8064 6190
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7104 5296 7156 5302
rect 7102 5264 7104 5273
rect 7156 5264 7158 5273
rect 7102 5199 7158 5208
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6472 4690 6500 4966
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 8220 4622 8248 5034
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 6012 3738 6040 4558
rect 7214 4380 7522 4389
rect 7214 4378 7220 4380
rect 7276 4378 7300 4380
rect 7356 4378 7380 4380
rect 7436 4378 7460 4380
rect 7516 4378 7522 4380
rect 7276 4326 7278 4378
rect 7458 4326 7460 4378
rect 7214 4324 7220 4326
rect 7276 4324 7300 4326
rect 7356 4324 7380 4326
rect 7436 4324 7460 4326
rect 7516 4324 7522 4326
rect 7214 4315 7522 4324
rect 8220 4282 8248 4558
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8220 4162 8248 4218
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 8128 4134 8248 4162
rect 7668 4049 7696 4082
rect 7932 4072 7984 4078
rect 7654 4040 7710 4049
rect 7932 4014 7984 4020
rect 7654 3975 7710 3984
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3738 7696 3878
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3896 2990 3924 3402
rect 4540 3194 4568 3402
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 5092 3126 5120 3402
rect 6932 3194 6960 3470
rect 7214 3292 7522 3301
rect 7214 3290 7220 3292
rect 7276 3290 7300 3292
rect 7356 3290 7380 3292
rect 7436 3290 7460 3292
rect 7516 3290 7522 3292
rect 7276 3238 7278 3290
rect 7458 3238 7460 3290
rect 7214 3236 7220 3238
rect 7276 3236 7300 3238
rect 7356 3236 7380 3238
rect 7436 3236 7460 3238
rect 7516 3236 7522 3238
rect 7214 3227 7522 3236
rect 7944 3194 7972 4014
rect 8128 3398 8156 4134
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8220 3738 8248 4014
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8312 3534 8340 8298
rect 8496 7818 8524 8366
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8588 7546 8616 8774
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8496 5302 8524 5510
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8588 5234 8616 5510
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 8680 3058 8708 4014
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8772 2650 8800 12038
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10742 9076 10950
rect 9232 10810 9260 11290
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9232 10062 9260 10746
rect 9508 10266 9536 12174
rect 9600 11354 9628 13126
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9876 12442 9904 12718
rect 9968 12646 9996 13670
rect 10214 13628 10522 13637
rect 10214 13626 10220 13628
rect 10276 13626 10300 13628
rect 10356 13626 10380 13628
rect 10436 13626 10460 13628
rect 10516 13626 10522 13628
rect 10276 13574 10278 13626
rect 10458 13574 10460 13626
rect 10214 13572 10220 13574
rect 10276 13572 10300 13574
rect 10356 13572 10380 13574
rect 10436 13572 10460 13574
rect 10516 13572 10522 13574
rect 10214 13563 10522 13572
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10520 12646 10548 13194
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9876 10810 9904 11018
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 8566 9352 9862
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 7410 8984 8230
rect 9324 7410 9352 8502
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9416 7206 9444 7754
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9048 5234 9076 5646
rect 9416 5522 9444 7142
rect 9508 5710 9536 9998
rect 9692 8974 9720 9998
rect 9784 9722 9812 10066
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9876 9382 9904 10746
rect 9968 9586 9996 12582
rect 10214 12540 10522 12549
rect 10214 12538 10220 12540
rect 10276 12538 10300 12540
rect 10356 12538 10380 12540
rect 10436 12538 10460 12540
rect 10516 12538 10522 12540
rect 10276 12486 10278 12538
rect 10458 12486 10460 12538
rect 10214 12484 10220 12486
rect 10276 12484 10300 12486
rect 10356 12484 10380 12486
rect 10436 12484 10460 12486
rect 10516 12484 10522 12486
rect 10214 12475 10522 12484
rect 10214 11452 10522 11461
rect 10214 11450 10220 11452
rect 10276 11450 10300 11452
rect 10356 11450 10380 11452
rect 10436 11450 10460 11452
rect 10516 11450 10522 11452
rect 10276 11398 10278 11450
rect 10458 11398 10460 11450
rect 10214 11396 10220 11398
rect 10276 11396 10300 11398
rect 10356 11396 10380 11398
rect 10436 11396 10460 11398
rect 10516 11396 10522 11398
rect 10214 11387 10522 11396
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 10606 10088 11154
rect 10612 10690 10640 13790
rect 10704 13462 10732 14010
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12238 10732 13126
rect 10796 12306 10824 13262
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12986 10916 13194
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10888 12442 10916 12922
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10980 11370 11008 15098
rect 11072 14278 11100 15438
rect 11164 14958 11192 15642
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11532 15450 11560 15506
rect 11532 15422 11744 15450
rect 11716 15366 11744 15422
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11716 15026 11744 15302
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11808 14958 11836 15642
rect 13096 15434 13124 16390
rect 13214 16348 13522 16357
rect 13214 16346 13220 16348
rect 13276 16346 13300 16348
rect 13356 16346 13380 16348
rect 13436 16346 13460 16348
rect 13516 16346 13522 16348
rect 13276 16294 13278 16346
rect 13458 16294 13460 16346
rect 13214 16292 13220 16294
rect 13276 16292 13300 16294
rect 13356 16292 13380 16294
rect 13436 16292 13460 16294
rect 13516 16292 13522 16294
rect 13214 16283 13522 16292
rect 13740 15706 13768 16730
rect 15488 16590 15516 18702
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 14384 16114 14412 16526
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14476 16182 14504 16390
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 12716 15428 12768 15434
rect 12716 15370 12768 15376
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12176 14618 12204 14758
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 11348 14414 11376 14554
rect 12268 14482 12296 14554
rect 12360 14482 12388 14758
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12348 14476 12400 14482
rect 12348 14418 12400 14424
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 12728 14346 12756 15370
rect 13214 15260 13522 15269
rect 13214 15258 13220 15260
rect 13276 15258 13300 15260
rect 13356 15258 13380 15260
rect 13436 15258 13460 15260
rect 13516 15258 13522 15260
rect 13276 15206 13278 15258
rect 13458 15206 13460 15258
rect 13214 15204 13220 15206
rect 13276 15204 13300 15206
rect 13356 15204 13380 15206
rect 13436 15204 13460 15206
rect 13516 15204 13522 15206
rect 13214 15195 13522 15204
rect 14108 15162 14136 15506
rect 14384 15162 14412 16050
rect 14752 15978 14780 16390
rect 14844 16250 14872 16390
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14752 15706 14780 15914
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14844 15502 14872 16186
rect 15028 16046 15056 16526
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15304 16250 15332 16458
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 15706 15424 15846
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 10888 11342 11008 11370
rect 11072 11354 11100 14214
rect 12728 14006 12756 14282
rect 13214 14172 13522 14181
rect 13214 14170 13220 14172
rect 13276 14170 13300 14172
rect 13356 14170 13380 14172
rect 13436 14170 13460 14172
rect 13516 14170 13522 14172
rect 13276 14118 13278 14170
rect 13458 14118 13460 14170
rect 13214 14116 13220 14118
rect 13276 14116 13300 14118
rect 13356 14116 13380 14118
rect 13436 14116 13460 14118
rect 13516 14116 13522 14118
rect 13214 14107 13522 14116
rect 14108 14074 14136 15098
rect 15488 15094 15516 15574
rect 15580 15502 15608 19450
rect 15936 19440 15988 19446
rect 15936 19382 15988 19388
rect 15948 18426 15976 19382
rect 16132 18766 16160 19722
rect 17788 19514 17816 20470
rect 17972 20262 18000 20810
rect 18156 20534 18184 21490
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17972 19514 18000 20198
rect 18156 20058 18184 20470
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 18156 19446 18184 19994
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 16214 19068 16522 19077
rect 16214 19066 16220 19068
rect 16276 19066 16300 19068
rect 16356 19066 16380 19068
rect 16436 19066 16460 19068
rect 16516 19066 16522 19068
rect 16276 19014 16278 19066
rect 16458 19014 16460 19066
rect 16214 19012 16220 19014
rect 16276 19012 16300 19014
rect 16356 19012 16380 19014
rect 16436 19012 16460 19014
rect 16516 19012 16522 19014
rect 16214 19003 16522 19012
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16132 18358 16160 18702
rect 16960 18426 16988 18906
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15672 17678 15700 18158
rect 16132 17882 16160 18294
rect 16960 18086 16988 18362
rect 17052 18358 17080 18566
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16214 17980 16522 17989
rect 16214 17978 16220 17980
rect 16276 17978 16300 17980
rect 16356 17978 16380 17980
rect 16436 17978 16460 17980
rect 16516 17978 16522 17980
rect 16276 17926 16278 17978
rect 16458 17926 16460 17978
rect 16214 17924 16220 17926
rect 16276 17924 16300 17926
rect 16356 17924 16380 17926
rect 16436 17924 16460 17926
rect 16516 17924 16522 17926
rect 16214 17915 16522 17924
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 16684 17610 16712 18022
rect 16960 17678 16988 18022
rect 17972 17882 18000 19110
rect 18248 18970 18276 21286
rect 18340 20466 18368 21286
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18340 20058 18368 20402
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18340 19446 18368 19994
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 18064 17746 18092 18226
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16868 17338 16896 17546
rect 18064 17338 18092 17682
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 16214 16892 16522 16901
rect 16214 16890 16220 16892
rect 16276 16890 16300 16892
rect 16356 16890 16380 16892
rect 16436 16890 16460 16892
rect 16516 16890 16522 16892
rect 16276 16838 16278 16890
rect 16458 16838 16460 16890
rect 16214 16836 16220 16838
rect 16276 16836 16300 16838
rect 16356 16836 16380 16838
rect 16436 16836 16460 16838
rect 16516 16836 16522 16838
rect 16214 16827 16522 16836
rect 16868 16794 16896 17274
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15672 15638 15700 16526
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15948 15706 15976 16186
rect 16040 16182 16068 16458
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15660 15632 15712 15638
rect 15660 15574 15712 15580
rect 16040 15570 16068 16118
rect 16214 15804 16522 15813
rect 16214 15802 16220 15804
rect 16276 15802 16300 15804
rect 16356 15802 16380 15804
rect 16436 15802 16460 15804
rect 16516 15802 16522 15804
rect 16276 15750 16278 15802
rect 16458 15750 16460 15802
rect 16214 15748 16220 15750
rect 16276 15748 16300 15750
rect 16356 15748 16380 15750
rect 16436 15748 16460 15750
rect 16516 15748 16522 15750
rect 16214 15739 16522 15748
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16684 15162 16712 15302
rect 17144 15162 17172 16594
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17316 15972 17368 15978
rect 17316 15914 17368 15920
rect 17328 15706 17356 15914
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17420 15706 17448 15846
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17788 15162 17816 15846
rect 17880 15434 17908 16390
rect 18156 16182 18184 18566
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18248 16182 18276 17478
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18340 16590 18368 16934
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18248 15722 18276 15982
rect 18248 15694 18368 15722
rect 18340 15638 18368 15694
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 14752 14550 14780 14962
rect 14740 14544 14792 14550
rect 14740 14486 14792 14492
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11440 12986 11468 13330
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11060 11348 11112 11354
rect 10888 11218 10916 11342
rect 11060 11290 11112 11296
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10888 10810 10916 11154
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10520 10662 10640 10690
rect 10520 10606 10548 10662
rect 10980 10606 11008 11086
rect 11164 10810 11192 12854
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11532 12442 11560 12718
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10060 9926 10088 10542
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 7750 9628 8230
rect 9692 7954 9720 8298
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9600 7478 9628 7686
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9600 6458 9628 7414
rect 9692 7410 9720 7890
rect 10152 7478 10180 10542
rect 10214 10364 10522 10373
rect 10214 10362 10220 10364
rect 10276 10362 10300 10364
rect 10356 10362 10380 10364
rect 10436 10362 10460 10364
rect 10516 10362 10522 10364
rect 10276 10310 10278 10362
rect 10458 10310 10460 10362
rect 10214 10308 10220 10310
rect 10276 10308 10300 10310
rect 10356 10308 10380 10310
rect 10436 10308 10460 10310
rect 10516 10308 10522 10310
rect 10214 10299 10522 10308
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9722 10364 9998
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10214 9276 10522 9285
rect 10214 9274 10220 9276
rect 10276 9274 10300 9276
rect 10356 9274 10380 9276
rect 10436 9274 10460 9276
rect 10516 9274 10522 9276
rect 10276 9222 10278 9274
rect 10458 9222 10460 9274
rect 10214 9220 10220 9222
rect 10276 9220 10300 9222
rect 10356 9220 10380 9222
rect 10436 9220 10460 9222
rect 10516 9220 10522 9222
rect 10214 9211 10522 9220
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10796 8634 10824 8842
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 8634 11100 8774
rect 11256 8634 11284 12174
rect 12452 11354 12480 12174
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11762 12572 12038
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12544 11354 12572 11698
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10742 11376 11154
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11532 10674 11560 11290
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10130 11560 10610
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11624 9994 11652 10950
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12176 10062 12204 10746
rect 12452 10130 12480 11290
rect 12728 10810 12756 13942
rect 14108 13394 14136 14010
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15488 13462 15516 13942
rect 15764 13870 15792 14962
rect 16214 14716 16522 14725
rect 16214 14714 16220 14716
rect 16276 14714 16300 14716
rect 16356 14714 16380 14716
rect 16436 14714 16460 14716
rect 16516 14714 16522 14716
rect 16276 14662 16278 14714
rect 16458 14662 16460 14714
rect 16214 14660 16220 14662
rect 16276 14660 16300 14662
rect 16356 14660 16380 14662
rect 16436 14660 16460 14662
rect 16516 14660 16522 14662
rect 16214 14651 16522 14660
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15856 13870 15884 14282
rect 16684 14278 16712 15098
rect 17880 14890 17908 15370
rect 18248 15094 18276 15438
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 17316 14884 17368 14890
rect 17316 14826 17368 14832
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 13214 13084 13522 13093
rect 13214 13082 13220 13084
rect 13276 13082 13300 13084
rect 13356 13082 13380 13084
rect 13436 13082 13460 13084
rect 13516 13082 13522 13084
rect 13276 13030 13278 13082
rect 13458 13030 13460 13082
rect 13214 13028 13220 13030
rect 13276 13028 13300 13030
rect 13356 13028 13380 13030
rect 13436 13028 13460 13030
rect 13516 13028 13522 13030
rect 13214 13019 13522 13028
rect 14108 12850 14136 13330
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14752 12986 14780 13194
rect 15488 12986 15516 13398
rect 15764 13326 15792 13806
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 13372 12442 13400 12786
rect 13924 12442 13952 12786
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13214 11996 13522 12005
rect 13214 11994 13220 11996
rect 13276 11994 13300 11996
rect 13356 11994 13380 11996
rect 13436 11994 13460 11996
rect 13516 11994 13522 11996
rect 13276 11942 13278 11994
rect 13458 11942 13460 11994
rect 13214 11940 13220 11942
rect 13276 11940 13300 11942
rect 13356 11940 13380 11942
rect 13436 11940 13460 11942
rect 13516 11940 13522 11942
rect 13214 11931 13522 11940
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13832 11150 13860 11766
rect 13924 11558 13952 12378
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14108 11762 14136 12310
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11830 14504 12038
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 14660 11150 14688 12786
rect 14752 12374 14780 12922
rect 15764 12850 15792 13262
rect 15856 12986 15884 13806
rect 15948 13734 15976 14214
rect 16304 14068 16356 14074
rect 16132 14028 16304 14056
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15948 13326 15976 13670
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 12986 15976 13262
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16040 12918 16068 13874
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15212 11898 15240 12310
rect 15580 12238 15608 12582
rect 16132 12434 16160 14028
rect 16304 14010 16356 14016
rect 16684 13870 16712 14214
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16214 13628 16522 13637
rect 16214 13626 16220 13628
rect 16276 13626 16300 13628
rect 16356 13626 16380 13628
rect 16436 13626 16460 13628
rect 16516 13626 16522 13628
rect 16276 13574 16278 13626
rect 16458 13574 16460 13626
rect 16214 13572 16220 13574
rect 16276 13572 16300 13574
rect 16356 13572 16380 13574
rect 16436 13572 16460 13574
rect 16516 13572 16522 13574
rect 16214 13563 16522 13572
rect 16684 13326 16712 13806
rect 16960 13462 16988 13874
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16214 12540 16522 12549
rect 16214 12538 16220 12540
rect 16276 12538 16300 12540
rect 16356 12538 16380 12540
rect 16436 12538 16460 12540
rect 16516 12538 16522 12540
rect 16276 12486 16278 12538
rect 16458 12486 16460 12538
rect 16214 12484 16220 12486
rect 16276 12484 16300 12486
rect 16356 12484 16380 12486
rect 16436 12484 16460 12486
rect 16516 12484 16522 12486
rect 16214 12475 16522 12484
rect 16684 12434 16712 13262
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16960 12434 16988 12582
rect 16132 12406 16344 12434
rect 16684 12406 16988 12434
rect 16316 12238 16344 12406
rect 16960 12306 16988 12406
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15856 11898 15884 12106
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16224 11898 16252 12038
rect 16408 11898 16436 12174
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11898 16712 12038
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 13214 10908 13522 10917
rect 13214 10906 13220 10908
rect 13276 10906 13300 10908
rect 13356 10906 13380 10908
rect 13436 10906 13460 10908
rect 13516 10906 13522 10908
rect 13276 10854 13278 10906
rect 13458 10854 13460 10906
rect 13214 10852 13220 10854
rect 13276 10852 13300 10854
rect 13356 10852 13380 10854
rect 13436 10852 13460 10854
rect 13516 10852 13522 10854
rect 13214 10843 13522 10852
rect 13832 10810 13860 11086
rect 15304 11014 15332 11766
rect 15580 11642 15608 11834
rect 16960 11830 16988 12242
rect 17236 12238 17264 12854
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17328 11830 17356 14826
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17420 12918 17448 13126
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 18064 12850 18092 13670
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17880 12434 17908 12582
rect 17788 12406 17908 12434
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 15488 11614 15608 11642
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 15028 10674 15056 10950
rect 15304 10742 15332 10950
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15488 10674 15516 11614
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11082 16160 11494
rect 16214 11452 16522 11461
rect 16214 11450 16220 11452
rect 16276 11450 16300 11452
rect 16356 11450 16380 11452
rect 16436 11450 16460 11452
rect 16516 11450 16522 11452
rect 16276 11398 16278 11450
rect 16458 11398 16460 11450
rect 16214 11396 16220 11398
rect 16276 11396 16300 11398
rect 16356 11396 16380 11398
rect 16436 11396 16460 11398
rect 16516 11396 16522 11398
rect 16214 11387 16522 11396
rect 16960 11218 16988 11766
rect 17788 11694 17816 12406
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16316 10810 16344 11018
rect 16960 10810 16988 11154
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 13214 9820 13522 9829
rect 13214 9818 13220 9820
rect 13276 9818 13300 9820
rect 13356 9818 13380 9820
rect 13436 9818 13460 9820
rect 13516 9818 13522 9820
rect 13276 9766 13278 9818
rect 13458 9766 13460 9818
rect 13214 9764 13220 9766
rect 13276 9764 13300 9766
rect 13356 9764 13380 9766
rect 13436 9764 13460 9766
rect 13516 9764 13522 9766
rect 13214 9755 13522 9764
rect 14384 9654 14412 9930
rect 15028 9722 15056 10610
rect 15488 10266 15516 10610
rect 16214 10364 16522 10373
rect 16214 10362 16220 10364
rect 16276 10362 16300 10364
rect 16356 10362 16380 10364
rect 16436 10362 16460 10364
rect 16516 10362 16522 10364
rect 16276 10310 16278 10362
rect 16458 10310 16460 10362
rect 16214 10308 16220 10310
rect 16276 10308 16300 10310
rect 16356 10308 16380 10310
rect 16436 10308 16460 10310
rect 16516 10308 16522 10310
rect 16214 10299 16522 10308
rect 16960 10266 16988 10746
rect 18156 10266 18184 14894
rect 18248 14074 18276 15030
rect 18616 14618 18644 21286
rect 18788 21140 18840 21146
rect 18788 21082 18840 21088
rect 18800 19854 18828 21082
rect 19214 20700 19522 20709
rect 19214 20698 19220 20700
rect 19276 20698 19300 20700
rect 19356 20698 19380 20700
rect 19436 20698 19460 20700
rect 19516 20698 19522 20700
rect 19276 20646 19278 20698
rect 19458 20646 19460 20698
rect 19214 20644 19220 20646
rect 19276 20644 19300 20646
rect 19356 20644 19380 20646
rect 19436 20644 19460 20646
rect 19516 20644 19522 20646
rect 19214 20635 19522 20644
rect 19616 20256 19668 20262
rect 19616 20198 19668 20204
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18800 19514 18828 19790
rect 19214 19612 19522 19621
rect 19214 19610 19220 19612
rect 19276 19610 19300 19612
rect 19356 19610 19380 19612
rect 19436 19610 19460 19612
rect 19516 19610 19522 19612
rect 19276 19558 19278 19610
rect 19458 19558 19460 19610
rect 19214 19556 19220 19558
rect 19276 19556 19300 19558
rect 19356 19556 19380 19558
rect 19436 19556 19460 19558
rect 19516 19556 19522 19558
rect 19214 19547 19522 19556
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 19628 19446 19656 20198
rect 19616 19440 19668 19446
rect 19668 19400 19748 19428
rect 19616 19382 19668 19388
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19214 18524 19522 18533
rect 19214 18522 19220 18524
rect 19276 18522 19300 18524
rect 19356 18522 19380 18524
rect 19436 18522 19460 18524
rect 19516 18522 19522 18524
rect 19276 18470 19278 18522
rect 19458 18470 19460 18522
rect 19214 18468 19220 18470
rect 19276 18468 19300 18470
rect 19356 18468 19380 18470
rect 19436 18468 19460 18470
rect 19516 18468 19522 18470
rect 19214 18459 19522 18468
rect 19628 18426 19656 18906
rect 19720 18766 19748 19400
rect 19800 19168 19852 19174
rect 19800 19110 19852 19116
rect 19812 18766 19840 19110
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19800 18760 19852 18766
rect 19800 18702 19852 18708
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19628 17678 19656 18362
rect 19720 17678 19748 18702
rect 19812 18358 19840 18702
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 19812 17746 19840 18294
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19708 17672 19760 17678
rect 19904 17626 19932 18702
rect 19708 17614 19760 17620
rect 19214 17436 19522 17445
rect 19214 17434 19220 17436
rect 19276 17434 19300 17436
rect 19356 17434 19380 17436
rect 19436 17434 19460 17436
rect 19516 17434 19522 17436
rect 19276 17382 19278 17434
rect 19458 17382 19460 17434
rect 19214 17380 19220 17382
rect 19276 17380 19300 17382
rect 19356 17380 19380 17382
rect 19436 17380 19460 17382
rect 19516 17380 19522 17382
rect 19214 17371 19522 17380
rect 19628 17270 19656 17614
rect 19812 17610 19932 17626
rect 19800 17604 19932 17610
rect 19852 17598 19932 17604
rect 19800 17546 19852 17552
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19812 16998 19840 17546
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 20272 16590 20300 21490
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 21185 20484 21286
rect 20442 21176 20498 21185
rect 20442 21111 20498 21120
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 16114 19012 16390
rect 19214 16348 19522 16357
rect 19214 16346 19220 16348
rect 19276 16346 19300 16348
rect 19356 16346 19380 16348
rect 19436 16346 19460 16348
rect 19516 16346 19522 16348
rect 19276 16294 19278 16346
rect 19458 16294 19460 16346
rect 19214 16292 19220 16294
rect 19276 16292 19300 16294
rect 19356 16292 19380 16294
rect 19436 16292 19460 16294
rect 19516 16292 19522 16294
rect 19214 16283 19522 16292
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 18696 15904 18748 15910
rect 18696 15846 18748 15852
rect 18708 15502 18736 15846
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18800 15162 18828 15438
rect 18892 15366 18920 15642
rect 18984 15502 19012 16050
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 19628 15366 19656 15846
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 18892 15026 18920 15302
rect 19214 15260 19522 15269
rect 19214 15258 19220 15260
rect 19276 15258 19300 15260
rect 19356 15258 19380 15260
rect 19436 15258 19460 15260
rect 19516 15258 19522 15260
rect 19276 15206 19278 15258
rect 19458 15206 19460 15258
rect 19214 15204 19220 15206
rect 19276 15204 19300 15206
rect 19356 15204 19380 15206
rect 19436 15204 19460 15206
rect 19516 15204 19522 15206
rect 19214 15195 19522 15204
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18892 14074 18920 14962
rect 19214 14172 19522 14181
rect 19214 14170 19220 14172
rect 19276 14170 19300 14172
rect 19356 14170 19380 14172
rect 19436 14170 19460 14172
rect 19516 14170 19522 14172
rect 19276 14118 19278 14170
rect 19458 14118 19460 14170
rect 19214 14116 19220 14118
rect 19276 14116 19300 14118
rect 19356 14116 19380 14118
rect 19436 14116 19460 14118
rect 19516 14116 19522 14118
rect 19214 14107 19522 14116
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 19628 14006 19656 15302
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 20272 13530 20300 15438
rect 20364 15094 20392 16050
rect 20442 15736 20498 15745
rect 20442 15671 20444 15680
rect 20496 15671 20498 15680
rect 20444 15642 20496 15648
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20260 13524 20312 13530
rect 20260 13466 20312 13472
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 18340 12918 18368 13194
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18340 12442 18368 12854
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18340 11762 18368 12038
rect 18524 11898 18552 12038
rect 18892 11898 18920 12378
rect 18984 12238 19012 12786
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 19076 11898 19104 13262
rect 19214 13084 19522 13093
rect 19214 13082 19220 13084
rect 19276 13082 19300 13084
rect 19356 13082 19380 13084
rect 19436 13082 19460 13084
rect 19516 13082 19522 13084
rect 19276 13030 19278 13082
rect 19458 13030 19460 13082
rect 19214 13028 19220 13030
rect 19276 13028 19300 13030
rect 19356 13028 19380 13030
rect 19436 13028 19460 13030
rect 19516 13028 19522 13030
rect 19214 13019 19522 13028
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19352 12306 19380 12922
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19214 11996 19522 12005
rect 19214 11994 19220 11996
rect 19276 11994 19300 11996
rect 19356 11994 19380 11996
rect 19436 11994 19460 11996
rect 19516 11994 19522 11996
rect 19276 11942 19278 11994
rect 19458 11942 19460 11994
rect 19214 11940 19220 11942
rect 19276 11940 19300 11942
rect 19356 11940 19380 11942
rect 19436 11940 19460 11942
rect 19516 11940 19522 11942
rect 19214 11931 19522 11940
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19628 11830 19656 12174
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18340 11558 18368 11698
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 10796 8378 10824 8434
rect 10796 8350 11100 8378
rect 10214 8188 10522 8197
rect 10214 8186 10220 8188
rect 10276 8186 10300 8188
rect 10356 8186 10380 8188
rect 10436 8186 10460 8188
rect 10516 8186 10522 8188
rect 10276 8134 10278 8186
rect 10458 8134 10460 8186
rect 10214 8132 10220 8134
rect 10276 8132 10300 8134
rect 10356 8132 10380 8134
rect 10436 8132 10460 8134
rect 10516 8132 10522 8134
rect 10214 8123 10522 8132
rect 11072 7818 11100 8350
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 8022 11376 8230
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 11624 7410 11652 8434
rect 11716 8090 11744 8434
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 12176 7954 12204 8774
rect 13214 8732 13522 8741
rect 13214 8730 13220 8732
rect 13276 8730 13300 8732
rect 13356 8730 13380 8732
rect 13436 8730 13460 8732
rect 13516 8730 13522 8732
rect 13276 8678 13278 8730
rect 13458 8678 13460 8730
rect 13214 8676 13220 8678
rect 13276 8676 13300 8678
rect 13356 8676 13380 8678
rect 13436 8676 13460 8678
rect 13516 8676 13522 8678
rect 13214 8667 13522 8676
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12452 7954 12480 8570
rect 13740 8498 13768 8842
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11808 7546 11836 7822
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 10214 7100 10522 7109
rect 10214 7098 10220 7100
rect 10276 7098 10300 7100
rect 10356 7098 10380 7100
rect 10436 7098 10460 7100
rect 10516 7098 10522 7100
rect 10276 7046 10278 7098
rect 10458 7046 10460 7098
rect 10214 7044 10220 7046
rect 10276 7044 10300 7046
rect 10356 7044 10380 7046
rect 10436 7044 10460 7046
rect 10516 7044 10522 7046
rect 10214 7035 10522 7044
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10214 6012 10522 6021
rect 10214 6010 10220 6012
rect 10276 6010 10300 6012
rect 10356 6010 10380 6012
rect 10436 6010 10460 6012
rect 10516 6010 10522 6012
rect 10276 5958 10278 6010
rect 10458 5958 10460 6010
rect 10214 5956 10220 5958
rect 10276 5956 10300 5958
rect 10356 5956 10380 5958
rect 10436 5956 10460 5958
rect 10516 5956 10522 5958
rect 10214 5947 10522 5956
rect 10704 5710 10732 6054
rect 11072 5914 11100 6190
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 9324 5494 9444 5522
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9048 4622 9076 5170
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 9140 4554 9168 4966
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9128 4548 9180 4554
rect 9128 4490 9180 4496
rect 9140 3466 9168 4490
rect 9232 3942 9260 4558
rect 9324 4146 9352 5494
rect 9508 5302 9536 5646
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 5302 9996 5510
rect 10060 5370 10088 5646
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9416 4622 9444 5170
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9508 4826 9536 4966
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9232 3466 9260 3878
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9324 3398 9352 4082
rect 9416 4078 9444 4558
rect 9692 4554 9720 5170
rect 10214 4924 10522 4933
rect 10214 4922 10220 4924
rect 10276 4922 10300 4924
rect 10356 4922 10380 4924
rect 10436 4922 10460 4924
rect 10516 4922 10522 4924
rect 10276 4870 10278 4922
rect 10458 4870 10460 4922
rect 10214 4868 10220 4870
rect 10276 4868 10300 4870
rect 10356 4868 10380 4870
rect 10436 4868 10460 4870
rect 10516 4868 10522 4870
rect 10214 4859 10522 4868
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9404 4072 9456 4078
rect 9692 4049 9720 4490
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9968 4146 9996 4422
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9404 4014 9456 4020
rect 9678 4040 9734 4049
rect 9416 3534 9444 4014
rect 9678 3975 9734 3984
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 9968 3738 9996 3878
rect 10214 3836 10522 3845
rect 10214 3834 10220 3836
rect 10276 3834 10300 3836
rect 10356 3834 10380 3836
rect 10436 3834 10460 3836
rect 10516 3834 10522 3836
rect 10276 3782 10278 3834
rect 10458 3782 10460 3834
rect 10214 3780 10220 3782
rect 10276 3780 10300 3782
rect 10356 3780 10380 3782
rect 10436 3780 10460 3782
rect 10516 3780 10522 3782
rect 10214 3771 10522 3780
rect 10612 3738 10640 3878
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9968 3398 9996 3674
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9324 3058 9352 3334
rect 10428 3194 10456 3538
rect 10704 3194 10732 3946
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 9692 2514 9720 2926
rect 11624 2922 11652 7346
rect 12452 5914 12480 7890
rect 13740 7818 13768 8434
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13832 8090 13860 8366
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 14108 7886 14136 8910
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13214 7644 13522 7653
rect 13214 7642 13220 7644
rect 13276 7642 13300 7644
rect 13356 7642 13380 7644
rect 13436 7642 13460 7644
rect 13516 7642 13522 7644
rect 13276 7590 13278 7642
rect 13458 7590 13460 7642
rect 13214 7588 13220 7590
rect 13276 7588 13300 7590
rect 13356 7588 13380 7590
rect 13436 7588 13460 7590
rect 13516 7588 13522 7590
rect 13214 7579 13522 7588
rect 13740 7206 13768 7754
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12820 6458 12848 6734
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 6458 12940 6598
rect 13214 6556 13522 6565
rect 13214 6554 13220 6556
rect 13276 6554 13300 6556
rect 13356 6554 13380 6556
rect 13436 6554 13460 6556
rect 13516 6554 13522 6556
rect 13276 6502 13278 6554
rect 13458 6502 13460 6554
rect 13214 6500 13220 6502
rect 13276 6500 13300 6502
rect 13356 6500 13380 6502
rect 13436 6500 13460 6502
rect 13516 6500 13522 6502
rect 13214 6491 13522 6500
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12636 5914 12664 6190
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12820 5846 12848 6394
rect 13740 6322 13768 7142
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 13004 5710 13032 6054
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 11716 5370 11744 5646
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 12176 5234 12204 5646
rect 12636 5574 12664 5646
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12544 5302 12572 5510
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12636 5234 12664 5510
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12176 4282 12204 5170
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3738 11928 3878
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11992 3618 12020 4014
rect 11900 3590 12112 3618
rect 11900 3398 11928 3590
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11808 3194 11836 3334
rect 11992 3194 12020 3470
rect 12084 3194 12112 3590
rect 12176 3380 12204 4218
rect 12636 4214 12664 5034
rect 13004 4622 13032 5646
rect 13096 5370 13124 5646
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13214 5468 13522 5477
rect 13214 5466 13220 5468
rect 13276 5466 13300 5468
rect 13356 5466 13380 5468
rect 13436 5466 13460 5468
rect 13516 5466 13522 5468
rect 13276 5414 13278 5466
rect 13458 5414 13460 5466
rect 13214 5412 13220 5414
rect 13276 5412 13300 5414
rect 13356 5412 13380 5414
rect 13436 5412 13460 5414
rect 13516 5412 13522 5414
rect 13214 5403 13522 5412
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13188 4826 13216 5102
rect 13740 5030 13768 5510
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13372 4622 13400 4966
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 13096 4146 13124 4558
rect 14200 4554 14228 9522
rect 14384 8974 14412 9590
rect 17972 9586 18000 9862
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 16214 9276 16522 9285
rect 16214 9274 16220 9276
rect 16276 9274 16300 9276
rect 16356 9274 16380 9276
rect 16436 9274 16460 9276
rect 16516 9274 16522 9276
rect 16276 9222 16278 9274
rect 16458 9222 16460 9274
rect 16214 9220 16220 9222
rect 16276 9220 16300 9222
rect 16356 9220 16380 9222
rect 16436 9220 16460 9222
rect 16516 9220 16522 9222
rect 16214 9211 16522 9220
rect 17420 9178 17448 9522
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15488 8566 15516 8774
rect 15764 8566 15792 8774
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15488 7886 15516 8502
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7410 15056 7686
rect 15764 7478 15792 8502
rect 16868 8294 16896 8842
rect 17604 8634 17632 8910
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17880 8498 17908 9046
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 16214 8188 16522 8197
rect 16214 8186 16220 8188
rect 16276 8186 16300 8188
rect 16356 8186 16380 8188
rect 16436 8186 16460 8188
rect 16516 8186 16522 8188
rect 16276 8134 16278 8186
rect 16458 8134 16460 8186
rect 16214 8132 16220 8134
rect 16276 8132 16300 8134
rect 16356 8132 16380 8134
rect 16436 8132 16460 8134
rect 16516 8132 16522 8134
rect 16214 8123 16522 8132
rect 16868 8090 16896 8230
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15028 6934 15056 7346
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 16132 6798 16160 7142
rect 16214 7100 16522 7109
rect 16214 7098 16220 7100
rect 16276 7098 16300 7100
rect 16356 7098 16380 7100
rect 16436 7098 16460 7100
rect 16516 7098 16522 7100
rect 16276 7046 16278 7098
rect 16458 7046 16460 7098
rect 16214 7044 16220 7046
rect 16276 7044 16300 7046
rect 16356 7044 16380 7046
rect 16436 7044 16460 7046
rect 16516 7044 16522 7046
rect 16214 7035 16522 7044
rect 17420 7002 17448 8230
rect 17880 8022 17908 8434
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17684 6996 17736 7002
rect 17684 6938 17736 6944
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16592 6118 16620 6666
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16214 6012 16522 6021
rect 16214 6010 16220 6012
rect 16276 6010 16300 6012
rect 16356 6010 16380 6012
rect 16436 6010 16460 6012
rect 16516 6010 16522 6012
rect 16276 5958 16278 6010
rect 16458 5958 16460 6010
rect 16214 5956 16220 5958
rect 16276 5956 16300 5958
rect 16356 5956 16380 5958
rect 16436 5956 16460 5958
rect 16516 5956 16522 5958
rect 16214 5947 16522 5956
rect 16592 5914 16620 6054
rect 16684 5914 16712 6802
rect 16948 6792 17000 6798
rect 17000 6740 17356 6746
rect 16948 6734 17356 6740
rect 16960 6730 17356 6734
rect 16960 6724 17368 6730
rect 16960 6718 17316 6724
rect 17316 6666 17368 6672
rect 17696 6662 17724 6938
rect 17972 6730 18000 9114
rect 18064 8294 18092 10066
rect 18248 9518 18276 10610
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18340 10062 18368 10406
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18340 9586 18368 9998
rect 18432 9722 18460 9998
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18340 8922 18368 9522
rect 18524 9382 18552 10678
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 9042 18552 9318
rect 18708 9178 18736 10066
rect 18892 9994 18920 11630
rect 19214 10908 19522 10917
rect 19214 10906 19220 10908
rect 19276 10906 19300 10908
rect 19356 10906 19380 10908
rect 19436 10906 19460 10908
rect 19516 10906 19522 10908
rect 19276 10854 19278 10906
rect 19458 10854 19460 10906
rect 19214 10852 19220 10854
rect 19276 10852 19300 10854
rect 19356 10852 19380 10854
rect 19436 10852 19460 10854
rect 19516 10852 19522 10854
rect 19214 10843 19522 10852
rect 20088 10674 20116 11834
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18892 9654 18920 9930
rect 19214 9820 19522 9829
rect 19214 9818 19220 9820
rect 19276 9818 19300 9820
rect 19356 9818 19380 9820
rect 19436 9818 19460 9820
rect 19516 9818 19522 9820
rect 19276 9766 19278 9818
rect 19458 9766 19460 9818
rect 19214 9764 19220 9766
rect 19276 9764 19300 9766
rect 19356 9764 19380 9766
rect 19436 9764 19460 9766
rect 19516 9764 19522 9766
rect 19214 9755 19522 9764
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 20088 9586 20116 10610
rect 20442 10296 20498 10305
rect 20442 10231 20498 10240
rect 20456 10130 20484 10231
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18340 8906 18552 8922
rect 18340 8900 18564 8906
rect 18340 8894 18512 8900
rect 18512 8842 18564 8848
rect 18800 8838 18828 9386
rect 18892 8838 18920 9454
rect 20088 9178 20116 9522
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18892 8498 18920 8774
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18156 8090 18184 8434
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18984 7886 19012 9046
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 19214 8732 19522 8741
rect 19214 8730 19220 8732
rect 19276 8730 19300 8732
rect 19356 8730 19380 8732
rect 19436 8730 19460 8732
rect 19516 8730 19522 8732
rect 19276 8678 19278 8730
rect 19458 8678 19460 8730
rect 19214 8676 19220 8678
rect 19276 8676 19300 8678
rect 19356 8676 19380 8678
rect 19436 8676 19460 8678
rect 19516 8676 19522 8678
rect 19214 8667 19522 8676
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19260 8090 19288 8502
rect 20364 8090 20392 8842
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18616 7546 18644 7754
rect 18984 7546 19012 7822
rect 19536 7750 19564 7890
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19214 7644 19522 7653
rect 19214 7642 19220 7644
rect 19276 7642 19300 7644
rect 19356 7642 19380 7644
rect 19436 7642 19460 7644
rect 19516 7642 19522 7644
rect 19276 7590 19278 7642
rect 19458 7590 19460 7642
rect 19214 7588 19220 7590
rect 19276 7588 19300 7590
rect 19356 7588 19380 7590
rect 19436 7588 19460 7590
rect 19516 7588 19522 7590
rect 19214 7579 19522 7588
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18420 7472 18472 7478
rect 18420 7414 18472 7420
rect 18432 7002 18460 7414
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17052 6458 17080 6598
rect 17696 6458 17724 6598
rect 18156 6458 18184 6734
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 17696 5642 17724 6394
rect 18432 6338 18460 6938
rect 19214 6556 19522 6565
rect 19214 6554 19220 6556
rect 19276 6554 19300 6556
rect 19356 6554 19380 6556
rect 19436 6554 19460 6556
rect 19516 6554 19522 6556
rect 19276 6502 19278 6554
rect 19458 6502 19460 6554
rect 19214 6500 19220 6502
rect 19276 6500 19300 6502
rect 19356 6500 19380 6502
rect 19436 6500 19460 6502
rect 19516 6500 19522 6502
rect 19214 6491 19522 6500
rect 18340 6322 18460 6338
rect 18328 6316 18460 6322
rect 18380 6310 18460 6316
rect 18328 6258 18380 6264
rect 19628 6118 19656 7822
rect 19720 7410 19748 7890
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 18156 5778 18184 6054
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 18156 5370 18184 5714
rect 19214 5468 19522 5477
rect 19214 5466 19220 5468
rect 19276 5466 19300 5468
rect 19356 5466 19380 5468
rect 19436 5466 19460 5468
rect 19516 5466 19522 5468
rect 19276 5414 19278 5466
rect 19458 5414 19460 5466
rect 19214 5412 19220 5414
rect 19276 5412 19300 5414
rect 19356 5412 19380 5414
rect 19436 5412 19460 5414
rect 19516 5412 19522 5414
rect 19214 5403 19522 5412
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 19628 5302 19656 6054
rect 19720 5370 19748 7346
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 14476 4758 14504 5238
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14752 4826 14780 5102
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 16214 4924 16522 4933
rect 16214 4922 16220 4924
rect 16276 4922 16300 4924
rect 16356 4922 16380 4924
rect 16436 4922 16460 4924
rect 16516 4922 16522 4924
rect 16276 4870 16278 4922
rect 16458 4870 16460 4922
rect 16214 4868 16220 4870
rect 16276 4868 16300 4870
rect 16356 4868 16380 4870
rect 16436 4868 16460 4870
rect 16516 4868 16522 4870
rect 16214 4859 16522 4868
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 13214 4380 13522 4389
rect 13214 4378 13220 4380
rect 13276 4378 13300 4380
rect 13356 4378 13380 4380
rect 13436 4378 13460 4380
rect 13516 4378 13522 4380
rect 13276 4326 13278 4378
rect 13458 4326 13460 4378
rect 13214 4324 13220 4326
rect 13276 4324 13300 4326
rect 13356 4324 13380 4326
rect 13436 4324 13460 4326
rect 13516 4324 13522 4326
rect 13214 4315 13522 4324
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12348 3392 12400 3398
rect 12176 3352 12348 3380
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12176 3074 12204 3352
rect 12348 3334 12400 3340
rect 11808 3058 12204 3074
rect 11796 3052 12204 3058
rect 11848 3046 12204 3052
rect 11796 2994 11848 3000
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 10214 2748 10522 2757
rect 10214 2746 10220 2748
rect 10276 2746 10300 2748
rect 10356 2746 10380 2748
rect 10436 2746 10460 2748
rect 10516 2746 10522 2748
rect 10276 2694 10278 2746
rect 10458 2694 10460 2746
rect 10214 2692 10220 2694
rect 10276 2692 10300 2694
rect 10356 2692 10380 2694
rect 10436 2692 10460 2694
rect 10516 2692 10522 2694
rect 10214 2683 10522 2692
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 12452 2446 12480 3878
rect 12544 3534 12572 3878
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 3126 12572 3334
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12544 2446 12572 3062
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12636 2650 12664 2926
rect 12728 2854 12756 3878
rect 13214 3292 13522 3301
rect 13214 3290 13220 3292
rect 13276 3290 13300 3292
rect 13356 3290 13380 3292
rect 13436 3290 13460 3292
rect 13516 3290 13522 3292
rect 13276 3238 13278 3290
rect 13458 3238 13460 3290
rect 13214 3236 13220 3238
rect 13276 3236 13300 3238
rect 13356 3236 13380 3238
rect 13436 3236 13460 3238
rect 13516 3236 13522 3238
rect 13214 3227 13522 3236
rect 14476 3176 14504 4694
rect 20272 4622 20300 4966
rect 20824 4865 20852 5170
rect 20810 4856 20866 4865
rect 20810 4791 20866 4800
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 19214 4380 19522 4389
rect 19214 4378 19220 4380
rect 19276 4378 19300 4380
rect 19356 4378 19380 4380
rect 19436 4378 19460 4380
rect 19516 4378 19522 4380
rect 19276 4326 19278 4378
rect 19458 4326 19460 4378
rect 19214 4324 19220 4326
rect 19276 4324 19300 4326
rect 19356 4324 19380 4326
rect 19436 4324 19460 4326
rect 19516 4324 19522 4326
rect 19214 4315 19522 4324
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 16214 3836 16522 3845
rect 16214 3834 16220 3836
rect 16276 3834 16300 3836
rect 16356 3834 16380 3836
rect 16436 3834 16460 3836
rect 16516 3834 16522 3836
rect 16276 3782 16278 3834
rect 16458 3782 16460 3834
rect 16214 3780 16220 3782
rect 16276 3780 16300 3782
rect 16356 3780 16380 3782
rect 16436 3780 16460 3782
rect 16516 3780 16522 3782
rect 16214 3771 16522 3780
rect 19214 3292 19522 3301
rect 19214 3290 19220 3292
rect 19276 3290 19300 3292
rect 19356 3290 19380 3292
rect 19436 3290 19460 3292
rect 19516 3290 19522 3292
rect 19276 3238 19278 3290
rect 19458 3238 19460 3290
rect 19214 3236 19220 3238
rect 19276 3236 19300 3238
rect 19356 3236 19380 3238
rect 19436 3236 19460 3238
rect 19516 3236 19522 3238
rect 19214 3227 19522 3236
rect 14556 3188 14608 3194
rect 14476 3148 14556 3176
rect 14556 3130 14608 3136
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 14200 2650 14228 2926
rect 14936 2774 14964 3062
rect 14936 2746 15240 2774
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 15212 2446 15240 2746
rect 16214 2748 16522 2757
rect 16214 2746 16220 2748
rect 16276 2746 16300 2748
rect 16356 2746 16380 2748
rect 16436 2746 16460 2748
rect 16516 2746 16522 2748
rect 16276 2694 16278 2746
rect 16458 2694 16460 2746
rect 16214 2692 16220 2694
rect 16276 2692 16300 2694
rect 16356 2692 16380 2694
rect 16436 2692 16460 2694
rect 16516 2692 16522 2694
rect 16214 2683 16522 2692
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 5276 1306 5304 2382
rect 7214 2204 7522 2213
rect 7214 2202 7220 2204
rect 7276 2202 7300 2204
rect 7356 2202 7380 2204
rect 7436 2202 7460 2204
rect 7516 2202 7522 2204
rect 7276 2150 7278 2202
rect 7458 2150 7460 2202
rect 7214 2148 7220 2150
rect 7276 2148 7300 2150
rect 7356 2148 7380 2150
rect 7436 2148 7460 2150
rect 7516 2148 7522 2150
rect 7214 2139 7522 2148
rect 10428 1306 10456 2382
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 13214 2204 13522 2213
rect 13214 2202 13220 2204
rect 13276 2202 13300 2204
rect 13356 2202 13380 2204
rect 13436 2202 13460 2204
rect 13516 2202 13522 2204
rect 13276 2150 13278 2202
rect 13458 2150 13460 2202
rect 13214 2148 13220 2150
rect 13276 2148 13300 2150
rect 13356 2148 13380 2150
rect 13436 2148 13460 2150
rect 13516 2148 13522 2150
rect 13214 2139 13522 2148
rect 5184 1278 5304 1306
rect 10336 1278 10456 1306
rect 5184 800 5212 1278
rect 10336 800 10364 1278
rect 15580 1170 15608 2314
rect 19214 2204 19522 2213
rect 19214 2202 19220 2204
rect 19276 2202 19300 2204
rect 19356 2202 19380 2204
rect 19436 2202 19460 2204
rect 19516 2202 19522 2204
rect 19276 2150 19278 2202
rect 19458 2150 19460 2202
rect 19214 2148 19220 2150
rect 19276 2148 19300 2150
rect 19356 2148 19380 2150
rect 19436 2148 19460 2150
rect 19516 2148 19522 2150
rect 19214 2139 19522 2148
rect 15488 1142 15608 1170
rect 15488 800 15516 1142
rect 20640 800 20668 4014
rect 18 0 74 800
rect 5170 0 5226 800
rect 10322 0 10378 800
rect 15474 0 15530 800
rect 20626 0 20682 800
<< via2 >>
rect 3146 21800 3202 21856
rect 938 16360 994 16416
rect 1398 10920 1454 10976
rect 7220 21786 7276 21788
rect 7300 21786 7356 21788
rect 7380 21786 7436 21788
rect 7460 21786 7516 21788
rect 7220 21734 7266 21786
rect 7266 21734 7276 21786
rect 7300 21734 7330 21786
rect 7330 21734 7342 21786
rect 7342 21734 7356 21786
rect 7380 21734 7394 21786
rect 7394 21734 7406 21786
rect 7406 21734 7436 21786
rect 7460 21734 7470 21786
rect 7470 21734 7516 21786
rect 7220 21732 7276 21734
rect 7300 21732 7356 21734
rect 7380 21732 7436 21734
rect 7460 21732 7516 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 13220 21786 13276 21788
rect 13300 21786 13356 21788
rect 13380 21786 13436 21788
rect 13460 21786 13516 21788
rect 13220 21734 13266 21786
rect 13266 21734 13276 21786
rect 13300 21734 13330 21786
rect 13330 21734 13342 21786
rect 13342 21734 13356 21786
rect 13380 21734 13394 21786
rect 13394 21734 13406 21786
rect 13406 21734 13436 21786
rect 13460 21734 13470 21786
rect 13470 21734 13516 21786
rect 13220 21732 13276 21734
rect 13300 21732 13356 21734
rect 13380 21732 13436 21734
rect 13460 21732 13516 21734
rect 19220 21786 19276 21788
rect 19300 21786 19356 21788
rect 19380 21786 19436 21788
rect 19460 21786 19516 21788
rect 19220 21734 19266 21786
rect 19266 21734 19276 21786
rect 19300 21734 19330 21786
rect 19330 21734 19342 21786
rect 19342 21734 19356 21786
rect 19380 21734 19394 21786
rect 19394 21734 19406 21786
rect 19406 21734 19436 21786
rect 19460 21734 19470 21786
rect 19470 21734 19516 21786
rect 19220 21732 19276 21734
rect 19300 21732 19356 21734
rect 19380 21732 19436 21734
rect 19460 21732 19516 21734
rect 10220 21242 10276 21244
rect 10300 21242 10356 21244
rect 10380 21242 10436 21244
rect 10460 21242 10516 21244
rect 10220 21190 10266 21242
rect 10266 21190 10276 21242
rect 10300 21190 10330 21242
rect 10330 21190 10342 21242
rect 10342 21190 10356 21242
rect 10380 21190 10394 21242
rect 10394 21190 10406 21242
rect 10406 21190 10436 21242
rect 10460 21190 10470 21242
rect 10470 21190 10516 21242
rect 10220 21188 10276 21190
rect 10300 21188 10356 21190
rect 10380 21188 10436 21190
rect 10460 21188 10516 21190
rect 16220 21242 16276 21244
rect 16300 21242 16356 21244
rect 16380 21242 16436 21244
rect 16460 21242 16516 21244
rect 16220 21190 16266 21242
rect 16266 21190 16276 21242
rect 16300 21190 16330 21242
rect 16330 21190 16342 21242
rect 16342 21190 16356 21242
rect 16380 21190 16394 21242
rect 16394 21190 16406 21242
rect 16406 21190 16436 21242
rect 16460 21190 16470 21242
rect 16470 21190 16516 21242
rect 16220 21188 16276 21190
rect 16300 21188 16356 21190
rect 16380 21188 16436 21190
rect 16460 21188 16516 21190
rect 7220 20698 7276 20700
rect 7300 20698 7356 20700
rect 7380 20698 7436 20700
rect 7460 20698 7516 20700
rect 7220 20646 7266 20698
rect 7266 20646 7276 20698
rect 7300 20646 7330 20698
rect 7330 20646 7342 20698
rect 7342 20646 7356 20698
rect 7380 20646 7394 20698
rect 7394 20646 7406 20698
rect 7406 20646 7436 20698
rect 7460 20646 7470 20698
rect 7470 20646 7516 20698
rect 7220 20644 7276 20646
rect 7300 20644 7356 20646
rect 7380 20644 7436 20646
rect 7460 20644 7516 20646
rect 7220 19610 7276 19612
rect 7300 19610 7356 19612
rect 7380 19610 7436 19612
rect 7460 19610 7516 19612
rect 7220 19558 7266 19610
rect 7266 19558 7276 19610
rect 7300 19558 7330 19610
rect 7330 19558 7342 19610
rect 7342 19558 7356 19610
rect 7380 19558 7394 19610
rect 7394 19558 7406 19610
rect 7406 19558 7436 19610
rect 7460 19558 7470 19610
rect 7470 19558 7516 19610
rect 7220 19556 7276 19558
rect 7300 19556 7356 19558
rect 7380 19556 7436 19558
rect 7460 19556 7516 19558
rect 10220 20154 10276 20156
rect 10300 20154 10356 20156
rect 10380 20154 10436 20156
rect 10460 20154 10516 20156
rect 10220 20102 10266 20154
rect 10266 20102 10276 20154
rect 10300 20102 10330 20154
rect 10330 20102 10342 20154
rect 10342 20102 10356 20154
rect 10380 20102 10394 20154
rect 10394 20102 10406 20154
rect 10406 20102 10436 20154
rect 10460 20102 10470 20154
rect 10470 20102 10516 20154
rect 10220 20100 10276 20102
rect 10300 20100 10356 20102
rect 10380 20100 10436 20102
rect 10460 20100 10516 20102
rect 7220 18522 7276 18524
rect 7300 18522 7356 18524
rect 7380 18522 7436 18524
rect 7460 18522 7516 18524
rect 7220 18470 7266 18522
rect 7266 18470 7276 18522
rect 7300 18470 7330 18522
rect 7330 18470 7342 18522
rect 7342 18470 7356 18522
rect 7380 18470 7394 18522
rect 7394 18470 7406 18522
rect 7406 18470 7436 18522
rect 7460 18470 7470 18522
rect 7470 18470 7516 18522
rect 7220 18468 7276 18470
rect 7300 18468 7356 18470
rect 7380 18468 7436 18470
rect 7460 18468 7516 18470
rect 13220 20698 13276 20700
rect 13300 20698 13356 20700
rect 13380 20698 13436 20700
rect 13460 20698 13516 20700
rect 13220 20646 13266 20698
rect 13266 20646 13276 20698
rect 13300 20646 13330 20698
rect 13330 20646 13342 20698
rect 13342 20646 13356 20698
rect 13380 20646 13394 20698
rect 13394 20646 13406 20698
rect 13406 20646 13436 20698
rect 13460 20646 13470 20698
rect 13470 20646 13516 20698
rect 13220 20644 13276 20646
rect 13300 20644 13356 20646
rect 13380 20644 13436 20646
rect 13460 20644 13516 20646
rect 13220 19610 13276 19612
rect 13300 19610 13356 19612
rect 13380 19610 13436 19612
rect 13460 19610 13516 19612
rect 13220 19558 13266 19610
rect 13266 19558 13276 19610
rect 13300 19558 13330 19610
rect 13330 19558 13342 19610
rect 13342 19558 13356 19610
rect 13380 19558 13394 19610
rect 13394 19558 13406 19610
rect 13406 19558 13436 19610
rect 13460 19558 13470 19610
rect 13470 19558 13516 19610
rect 13220 19556 13276 19558
rect 13300 19556 13356 19558
rect 13380 19556 13436 19558
rect 13460 19556 13516 19558
rect 10220 19066 10276 19068
rect 10300 19066 10356 19068
rect 10380 19066 10436 19068
rect 10460 19066 10516 19068
rect 10220 19014 10266 19066
rect 10266 19014 10276 19066
rect 10300 19014 10330 19066
rect 10330 19014 10342 19066
rect 10342 19014 10356 19066
rect 10380 19014 10394 19066
rect 10394 19014 10406 19066
rect 10406 19014 10436 19066
rect 10460 19014 10470 19066
rect 10470 19014 10516 19066
rect 10220 19012 10276 19014
rect 10300 19012 10356 19014
rect 10380 19012 10436 19014
rect 10460 19012 10516 19014
rect 13220 18522 13276 18524
rect 13300 18522 13356 18524
rect 13380 18522 13436 18524
rect 13460 18522 13516 18524
rect 13220 18470 13266 18522
rect 13266 18470 13276 18522
rect 13300 18470 13330 18522
rect 13330 18470 13342 18522
rect 13342 18470 13356 18522
rect 13380 18470 13394 18522
rect 13394 18470 13406 18522
rect 13406 18470 13436 18522
rect 13460 18470 13470 18522
rect 13470 18470 13516 18522
rect 13220 18468 13276 18470
rect 13300 18468 13356 18470
rect 13380 18468 13436 18470
rect 13460 18468 13516 18470
rect 7220 17434 7276 17436
rect 7300 17434 7356 17436
rect 7380 17434 7436 17436
rect 7460 17434 7516 17436
rect 7220 17382 7266 17434
rect 7266 17382 7276 17434
rect 7300 17382 7330 17434
rect 7330 17382 7342 17434
rect 7342 17382 7356 17434
rect 7380 17382 7394 17434
rect 7394 17382 7406 17434
rect 7406 17382 7436 17434
rect 7460 17382 7470 17434
rect 7470 17382 7516 17434
rect 7220 17380 7276 17382
rect 7300 17380 7356 17382
rect 7380 17380 7436 17382
rect 7460 17380 7516 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 10220 17978 10276 17980
rect 10300 17978 10356 17980
rect 10380 17978 10436 17980
rect 10460 17978 10516 17980
rect 10220 17926 10266 17978
rect 10266 17926 10276 17978
rect 10300 17926 10330 17978
rect 10330 17926 10342 17978
rect 10342 17926 10356 17978
rect 10380 17926 10394 17978
rect 10394 17926 10406 17978
rect 10406 17926 10436 17978
rect 10460 17926 10470 17978
rect 10470 17926 10516 17978
rect 10220 17924 10276 17926
rect 10300 17924 10356 17926
rect 10380 17924 10436 17926
rect 10460 17924 10516 17926
rect 13220 17434 13276 17436
rect 13300 17434 13356 17436
rect 13380 17434 13436 17436
rect 13460 17434 13516 17436
rect 13220 17382 13266 17434
rect 13266 17382 13276 17434
rect 13300 17382 13330 17434
rect 13330 17382 13342 17434
rect 13342 17382 13356 17434
rect 13380 17382 13394 17434
rect 13394 17382 13406 17434
rect 13406 17382 13436 17434
rect 13460 17382 13470 17434
rect 13470 17382 13516 17434
rect 13220 17380 13276 17382
rect 13300 17380 13356 17382
rect 13380 17380 13436 17382
rect 13460 17380 13516 17382
rect 7220 16346 7276 16348
rect 7300 16346 7356 16348
rect 7380 16346 7436 16348
rect 7460 16346 7516 16348
rect 7220 16294 7266 16346
rect 7266 16294 7276 16346
rect 7300 16294 7330 16346
rect 7330 16294 7342 16346
rect 7342 16294 7356 16346
rect 7380 16294 7394 16346
rect 7394 16294 7406 16346
rect 7406 16294 7436 16346
rect 7460 16294 7470 16346
rect 7470 16294 7516 16346
rect 7220 16292 7276 16294
rect 7300 16292 7356 16294
rect 7380 16292 7436 16294
rect 7460 16292 7516 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 7220 15258 7276 15260
rect 7300 15258 7356 15260
rect 7380 15258 7436 15260
rect 7460 15258 7516 15260
rect 7220 15206 7266 15258
rect 7266 15206 7276 15258
rect 7300 15206 7330 15258
rect 7330 15206 7342 15258
rect 7342 15206 7356 15258
rect 7380 15206 7394 15258
rect 7394 15206 7406 15258
rect 7406 15206 7436 15258
rect 7460 15206 7470 15258
rect 7470 15206 7516 15258
rect 7220 15204 7276 15206
rect 7300 15204 7356 15206
rect 7380 15204 7436 15206
rect 7460 15204 7516 15206
rect 7220 14170 7276 14172
rect 7300 14170 7356 14172
rect 7380 14170 7436 14172
rect 7460 14170 7516 14172
rect 7220 14118 7266 14170
rect 7266 14118 7276 14170
rect 7300 14118 7330 14170
rect 7330 14118 7342 14170
rect 7342 14118 7356 14170
rect 7380 14118 7394 14170
rect 7394 14118 7406 14170
rect 7406 14118 7436 14170
rect 7460 14118 7470 14170
rect 7470 14118 7516 14170
rect 7220 14116 7276 14118
rect 7300 14116 7356 14118
rect 7380 14116 7436 14118
rect 7460 14116 7516 14118
rect 1398 5480 1454 5536
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 7220 13082 7276 13084
rect 7300 13082 7356 13084
rect 7380 13082 7436 13084
rect 7460 13082 7516 13084
rect 7220 13030 7266 13082
rect 7266 13030 7276 13082
rect 7300 13030 7330 13082
rect 7330 13030 7342 13082
rect 7342 13030 7356 13082
rect 7380 13030 7394 13082
rect 7394 13030 7406 13082
rect 7406 13030 7436 13082
rect 7460 13030 7470 13082
rect 7470 13030 7516 13082
rect 7220 13028 7276 13030
rect 7300 13028 7356 13030
rect 7380 13028 7436 13030
rect 7460 13028 7516 13030
rect 7220 11994 7276 11996
rect 7300 11994 7356 11996
rect 7380 11994 7436 11996
rect 7460 11994 7516 11996
rect 7220 11942 7266 11994
rect 7266 11942 7276 11994
rect 7300 11942 7330 11994
rect 7330 11942 7342 11994
rect 7342 11942 7356 11994
rect 7380 11942 7394 11994
rect 7394 11942 7406 11994
rect 7406 11942 7436 11994
rect 7460 11942 7470 11994
rect 7470 11942 7516 11994
rect 7220 11940 7276 11942
rect 7300 11940 7356 11942
rect 7380 11940 7436 11942
rect 7460 11940 7516 11942
rect 7220 10906 7276 10908
rect 7300 10906 7356 10908
rect 7380 10906 7436 10908
rect 7460 10906 7516 10908
rect 7220 10854 7266 10906
rect 7266 10854 7276 10906
rect 7300 10854 7330 10906
rect 7330 10854 7342 10906
rect 7342 10854 7356 10906
rect 7380 10854 7394 10906
rect 7394 10854 7406 10906
rect 7406 10854 7436 10906
rect 7460 10854 7470 10906
rect 7470 10854 7516 10906
rect 7220 10852 7276 10854
rect 7300 10852 7356 10854
rect 7380 10852 7436 10854
rect 7460 10852 7516 10854
rect 7220 9818 7276 9820
rect 7300 9818 7356 9820
rect 7380 9818 7436 9820
rect 7460 9818 7516 9820
rect 7220 9766 7266 9818
rect 7266 9766 7276 9818
rect 7300 9766 7330 9818
rect 7330 9766 7342 9818
rect 7342 9766 7356 9818
rect 7380 9766 7394 9818
rect 7394 9766 7406 9818
rect 7406 9766 7436 9818
rect 7460 9766 7470 9818
rect 7470 9766 7516 9818
rect 7220 9764 7276 9766
rect 7300 9764 7356 9766
rect 7380 9764 7436 9766
rect 7460 9764 7516 9766
rect 7220 8730 7276 8732
rect 7300 8730 7356 8732
rect 7380 8730 7436 8732
rect 7460 8730 7516 8732
rect 7220 8678 7266 8730
rect 7266 8678 7276 8730
rect 7300 8678 7330 8730
rect 7330 8678 7342 8730
rect 7342 8678 7356 8730
rect 7380 8678 7394 8730
rect 7394 8678 7406 8730
rect 7406 8678 7436 8730
rect 7460 8678 7470 8730
rect 7470 8678 7516 8730
rect 7220 8676 7276 8678
rect 7300 8676 7356 8678
rect 7380 8676 7436 8678
rect 7460 8676 7516 8678
rect 10220 16890 10276 16892
rect 10300 16890 10356 16892
rect 10380 16890 10436 16892
rect 10460 16890 10516 16892
rect 10220 16838 10266 16890
rect 10266 16838 10276 16890
rect 10300 16838 10330 16890
rect 10330 16838 10342 16890
rect 10342 16838 10356 16890
rect 10380 16838 10394 16890
rect 10394 16838 10406 16890
rect 10406 16838 10436 16890
rect 10460 16838 10470 16890
rect 10470 16838 10516 16890
rect 10220 16836 10276 16838
rect 10300 16836 10356 16838
rect 10380 16836 10436 16838
rect 10460 16836 10516 16838
rect 10220 15802 10276 15804
rect 10300 15802 10356 15804
rect 10380 15802 10436 15804
rect 10460 15802 10516 15804
rect 10220 15750 10266 15802
rect 10266 15750 10276 15802
rect 10300 15750 10330 15802
rect 10330 15750 10342 15802
rect 10342 15750 10356 15802
rect 10380 15750 10394 15802
rect 10394 15750 10406 15802
rect 10406 15750 10436 15802
rect 10460 15750 10470 15802
rect 10470 15750 10516 15802
rect 10220 15748 10276 15750
rect 10300 15748 10356 15750
rect 10380 15748 10436 15750
rect 10460 15748 10516 15750
rect 16220 20154 16276 20156
rect 16300 20154 16356 20156
rect 16380 20154 16436 20156
rect 16460 20154 16516 20156
rect 16220 20102 16266 20154
rect 16266 20102 16276 20154
rect 16300 20102 16330 20154
rect 16330 20102 16342 20154
rect 16342 20102 16356 20154
rect 16380 20102 16394 20154
rect 16394 20102 16406 20154
rect 16406 20102 16436 20154
rect 16460 20102 16470 20154
rect 16470 20102 16516 20154
rect 16220 20100 16276 20102
rect 16300 20100 16356 20102
rect 16380 20100 16436 20102
rect 16460 20100 16516 20102
rect 10220 14714 10276 14716
rect 10300 14714 10356 14716
rect 10380 14714 10436 14716
rect 10460 14714 10516 14716
rect 10220 14662 10266 14714
rect 10266 14662 10276 14714
rect 10300 14662 10330 14714
rect 10330 14662 10342 14714
rect 10342 14662 10356 14714
rect 10380 14662 10394 14714
rect 10394 14662 10406 14714
rect 10406 14662 10436 14714
rect 10460 14662 10470 14714
rect 10470 14662 10516 14714
rect 10220 14660 10276 14662
rect 10300 14660 10356 14662
rect 10380 14660 10436 14662
rect 10460 14660 10516 14662
rect 7220 7642 7276 7644
rect 7300 7642 7356 7644
rect 7380 7642 7436 7644
rect 7460 7642 7516 7644
rect 7220 7590 7266 7642
rect 7266 7590 7276 7642
rect 7300 7590 7330 7642
rect 7330 7590 7342 7642
rect 7342 7590 7356 7642
rect 7380 7590 7394 7642
rect 7394 7590 7406 7642
rect 7406 7590 7436 7642
rect 7460 7590 7470 7642
rect 7470 7590 7516 7642
rect 7220 7588 7276 7590
rect 7300 7588 7356 7590
rect 7380 7588 7436 7590
rect 7460 7588 7516 7590
rect 7220 6554 7276 6556
rect 7300 6554 7356 6556
rect 7380 6554 7436 6556
rect 7460 6554 7516 6556
rect 7220 6502 7266 6554
rect 7266 6502 7276 6554
rect 7300 6502 7330 6554
rect 7330 6502 7342 6554
rect 7342 6502 7356 6554
rect 7380 6502 7394 6554
rect 7394 6502 7406 6554
rect 7406 6502 7436 6554
rect 7460 6502 7470 6554
rect 7470 6502 7516 6554
rect 7220 6500 7276 6502
rect 7300 6500 7356 6502
rect 7380 6500 7436 6502
rect 7460 6500 7516 6502
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 6274 5244 6276 5264
rect 6276 5244 6328 5264
rect 6328 5244 6330 5264
rect 6274 5208 6330 5244
rect 7220 5466 7276 5468
rect 7300 5466 7356 5468
rect 7380 5466 7436 5468
rect 7460 5466 7516 5468
rect 7220 5414 7266 5466
rect 7266 5414 7276 5466
rect 7300 5414 7330 5466
rect 7330 5414 7342 5466
rect 7342 5414 7356 5466
rect 7380 5414 7394 5466
rect 7394 5414 7406 5466
rect 7406 5414 7436 5466
rect 7460 5414 7470 5466
rect 7470 5414 7516 5466
rect 7220 5412 7276 5414
rect 7300 5412 7356 5414
rect 7380 5412 7436 5414
rect 7460 5412 7516 5414
rect 7102 5244 7104 5264
rect 7104 5244 7156 5264
rect 7156 5244 7158 5264
rect 7102 5208 7158 5244
rect 7220 4378 7276 4380
rect 7300 4378 7356 4380
rect 7380 4378 7436 4380
rect 7460 4378 7516 4380
rect 7220 4326 7266 4378
rect 7266 4326 7276 4378
rect 7300 4326 7330 4378
rect 7330 4326 7342 4378
rect 7342 4326 7356 4378
rect 7380 4326 7394 4378
rect 7394 4326 7406 4378
rect 7406 4326 7436 4378
rect 7460 4326 7470 4378
rect 7470 4326 7516 4378
rect 7220 4324 7276 4326
rect 7300 4324 7356 4326
rect 7380 4324 7436 4326
rect 7460 4324 7516 4326
rect 7654 3984 7710 4040
rect 7220 3290 7276 3292
rect 7300 3290 7356 3292
rect 7380 3290 7436 3292
rect 7460 3290 7516 3292
rect 7220 3238 7266 3290
rect 7266 3238 7276 3290
rect 7300 3238 7330 3290
rect 7330 3238 7342 3290
rect 7342 3238 7356 3290
rect 7380 3238 7394 3290
rect 7394 3238 7406 3290
rect 7406 3238 7436 3290
rect 7460 3238 7470 3290
rect 7470 3238 7516 3290
rect 7220 3236 7276 3238
rect 7300 3236 7356 3238
rect 7380 3236 7436 3238
rect 7460 3236 7516 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10220 13626 10276 13628
rect 10300 13626 10356 13628
rect 10380 13626 10436 13628
rect 10460 13626 10516 13628
rect 10220 13574 10266 13626
rect 10266 13574 10276 13626
rect 10300 13574 10330 13626
rect 10330 13574 10342 13626
rect 10342 13574 10356 13626
rect 10380 13574 10394 13626
rect 10394 13574 10406 13626
rect 10406 13574 10436 13626
rect 10460 13574 10470 13626
rect 10470 13574 10516 13626
rect 10220 13572 10276 13574
rect 10300 13572 10356 13574
rect 10380 13572 10436 13574
rect 10460 13572 10516 13574
rect 10220 12538 10276 12540
rect 10300 12538 10356 12540
rect 10380 12538 10436 12540
rect 10460 12538 10516 12540
rect 10220 12486 10266 12538
rect 10266 12486 10276 12538
rect 10300 12486 10330 12538
rect 10330 12486 10342 12538
rect 10342 12486 10356 12538
rect 10380 12486 10394 12538
rect 10394 12486 10406 12538
rect 10406 12486 10436 12538
rect 10460 12486 10470 12538
rect 10470 12486 10516 12538
rect 10220 12484 10276 12486
rect 10300 12484 10356 12486
rect 10380 12484 10436 12486
rect 10460 12484 10516 12486
rect 10220 11450 10276 11452
rect 10300 11450 10356 11452
rect 10380 11450 10436 11452
rect 10460 11450 10516 11452
rect 10220 11398 10266 11450
rect 10266 11398 10276 11450
rect 10300 11398 10330 11450
rect 10330 11398 10342 11450
rect 10342 11398 10356 11450
rect 10380 11398 10394 11450
rect 10394 11398 10406 11450
rect 10406 11398 10436 11450
rect 10460 11398 10470 11450
rect 10470 11398 10516 11450
rect 10220 11396 10276 11398
rect 10300 11396 10356 11398
rect 10380 11396 10436 11398
rect 10460 11396 10516 11398
rect 13220 16346 13276 16348
rect 13300 16346 13356 16348
rect 13380 16346 13436 16348
rect 13460 16346 13516 16348
rect 13220 16294 13266 16346
rect 13266 16294 13276 16346
rect 13300 16294 13330 16346
rect 13330 16294 13342 16346
rect 13342 16294 13356 16346
rect 13380 16294 13394 16346
rect 13394 16294 13406 16346
rect 13406 16294 13436 16346
rect 13460 16294 13470 16346
rect 13470 16294 13516 16346
rect 13220 16292 13276 16294
rect 13300 16292 13356 16294
rect 13380 16292 13436 16294
rect 13460 16292 13516 16294
rect 13220 15258 13276 15260
rect 13300 15258 13356 15260
rect 13380 15258 13436 15260
rect 13460 15258 13516 15260
rect 13220 15206 13266 15258
rect 13266 15206 13276 15258
rect 13300 15206 13330 15258
rect 13330 15206 13342 15258
rect 13342 15206 13356 15258
rect 13380 15206 13394 15258
rect 13394 15206 13406 15258
rect 13406 15206 13436 15258
rect 13460 15206 13470 15258
rect 13470 15206 13516 15258
rect 13220 15204 13276 15206
rect 13300 15204 13356 15206
rect 13380 15204 13436 15206
rect 13460 15204 13516 15206
rect 13220 14170 13276 14172
rect 13300 14170 13356 14172
rect 13380 14170 13436 14172
rect 13460 14170 13516 14172
rect 13220 14118 13266 14170
rect 13266 14118 13276 14170
rect 13300 14118 13330 14170
rect 13330 14118 13342 14170
rect 13342 14118 13356 14170
rect 13380 14118 13394 14170
rect 13394 14118 13406 14170
rect 13406 14118 13436 14170
rect 13460 14118 13470 14170
rect 13470 14118 13516 14170
rect 13220 14116 13276 14118
rect 13300 14116 13356 14118
rect 13380 14116 13436 14118
rect 13460 14116 13516 14118
rect 16220 19066 16276 19068
rect 16300 19066 16356 19068
rect 16380 19066 16436 19068
rect 16460 19066 16516 19068
rect 16220 19014 16266 19066
rect 16266 19014 16276 19066
rect 16300 19014 16330 19066
rect 16330 19014 16342 19066
rect 16342 19014 16356 19066
rect 16380 19014 16394 19066
rect 16394 19014 16406 19066
rect 16406 19014 16436 19066
rect 16460 19014 16470 19066
rect 16470 19014 16516 19066
rect 16220 19012 16276 19014
rect 16300 19012 16356 19014
rect 16380 19012 16436 19014
rect 16460 19012 16516 19014
rect 16220 17978 16276 17980
rect 16300 17978 16356 17980
rect 16380 17978 16436 17980
rect 16460 17978 16516 17980
rect 16220 17926 16266 17978
rect 16266 17926 16276 17978
rect 16300 17926 16330 17978
rect 16330 17926 16342 17978
rect 16342 17926 16356 17978
rect 16380 17926 16394 17978
rect 16394 17926 16406 17978
rect 16406 17926 16436 17978
rect 16460 17926 16470 17978
rect 16470 17926 16516 17978
rect 16220 17924 16276 17926
rect 16300 17924 16356 17926
rect 16380 17924 16436 17926
rect 16460 17924 16516 17926
rect 16220 16890 16276 16892
rect 16300 16890 16356 16892
rect 16380 16890 16436 16892
rect 16460 16890 16516 16892
rect 16220 16838 16266 16890
rect 16266 16838 16276 16890
rect 16300 16838 16330 16890
rect 16330 16838 16342 16890
rect 16342 16838 16356 16890
rect 16380 16838 16394 16890
rect 16394 16838 16406 16890
rect 16406 16838 16436 16890
rect 16460 16838 16470 16890
rect 16470 16838 16516 16890
rect 16220 16836 16276 16838
rect 16300 16836 16356 16838
rect 16380 16836 16436 16838
rect 16460 16836 16516 16838
rect 16220 15802 16276 15804
rect 16300 15802 16356 15804
rect 16380 15802 16436 15804
rect 16460 15802 16516 15804
rect 16220 15750 16266 15802
rect 16266 15750 16276 15802
rect 16300 15750 16330 15802
rect 16330 15750 16342 15802
rect 16342 15750 16356 15802
rect 16380 15750 16394 15802
rect 16394 15750 16406 15802
rect 16406 15750 16436 15802
rect 16460 15750 16470 15802
rect 16470 15750 16516 15802
rect 16220 15748 16276 15750
rect 16300 15748 16356 15750
rect 16380 15748 16436 15750
rect 16460 15748 16516 15750
rect 10220 10362 10276 10364
rect 10300 10362 10356 10364
rect 10380 10362 10436 10364
rect 10460 10362 10516 10364
rect 10220 10310 10266 10362
rect 10266 10310 10276 10362
rect 10300 10310 10330 10362
rect 10330 10310 10342 10362
rect 10342 10310 10356 10362
rect 10380 10310 10394 10362
rect 10394 10310 10406 10362
rect 10406 10310 10436 10362
rect 10460 10310 10470 10362
rect 10470 10310 10516 10362
rect 10220 10308 10276 10310
rect 10300 10308 10356 10310
rect 10380 10308 10436 10310
rect 10460 10308 10516 10310
rect 10220 9274 10276 9276
rect 10300 9274 10356 9276
rect 10380 9274 10436 9276
rect 10460 9274 10516 9276
rect 10220 9222 10266 9274
rect 10266 9222 10276 9274
rect 10300 9222 10330 9274
rect 10330 9222 10342 9274
rect 10342 9222 10356 9274
rect 10380 9222 10394 9274
rect 10394 9222 10406 9274
rect 10406 9222 10436 9274
rect 10460 9222 10470 9274
rect 10470 9222 10516 9274
rect 10220 9220 10276 9222
rect 10300 9220 10356 9222
rect 10380 9220 10436 9222
rect 10460 9220 10516 9222
rect 16220 14714 16276 14716
rect 16300 14714 16356 14716
rect 16380 14714 16436 14716
rect 16460 14714 16516 14716
rect 16220 14662 16266 14714
rect 16266 14662 16276 14714
rect 16300 14662 16330 14714
rect 16330 14662 16342 14714
rect 16342 14662 16356 14714
rect 16380 14662 16394 14714
rect 16394 14662 16406 14714
rect 16406 14662 16436 14714
rect 16460 14662 16470 14714
rect 16470 14662 16516 14714
rect 16220 14660 16276 14662
rect 16300 14660 16356 14662
rect 16380 14660 16436 14662
rect 16460 14660 16516 14662
rect 13220 13082 13276 13084
rect 13300 13082 13356 13084
rect 13380 13082 13436 13084
rect 13460 13082 13516 13084
rect 13220 13030 13266 13082
rect 13266 13030 13276 13082
rect 13300 13030 13330 13082
rect 13330 13030 13342 13082
rect 13342 13030 13356 13082
rect 13380 13030 13394 13082
rect 13394 13030 13406 13082
rect 13406 13030 13436 13082
rect 13460 13030 13470 13082
rect 13470 13030 13516 13082
rect 13220 13028 13276 13030
rect 13300 13028 13356 13030
rect 13380 13028 13436 13030
rect 13460 13028 13516 13030
rect 13220 11994 13276 11996
rect 13300 11994 13356 11996
rect 13380 11994 13436 11996
rect 13460 11994 13516 11996
rect 13220 11942 13266 11994
rect 13266 11942 13276 11994
rect 13300 11942 13330 11994
rect 13330 11942 13342 11994
rect 13342 11942 13356 11994
rect 13380 11942 13394 11994
rect 13394 11942 13406 11994
rect 13406 11942 13436 11994
rect 13460 11942 13470 11994
rect 13470 11942 13516 11994
rect 13220 11940 13276 11942
rect 13300 11940 13356 11942
rect 13380 11940 13436 11942
rect 13460 11940 13516 11942
rect 16220 13626 16276 13628
rect 16300 13626 16356 13628
rect 16380 13626 16436 13628
rect 16460 13626 16516 13628
rect 16220 13574 16266 13626
rect 16266 13574 16276 13626
rect 16300 13574 16330 13626
rect 16330 13574 16342 13626
rect 16342 13574 16356 13626
rect 16380 13574 16394 13626
rect 16394 13574 16406 13626
rect 16406 13574 16436 13626
rect 16460 13574 16470 13626
rect 16470 13574 16516 13626
rect 16220 13572 16276 13574
rect 16300 13572 16356 13574
rect 16380 13572 16436 13574
rect 16460 13572 16516 13574
rect 16220 12538 16276 12540
rect 16300 12538 16356 12540
rect 16380 12538 16436 12540
rect 16460 12538 16516 12540
rect 16220 12486 16266 12538
rect 16266 12486 16276 12538
rect 16300 12486 16330 12538
rect 16330 12486 16342 12538
rect 16342 12486 16356 12538
rect 16380 12486 16394 12538
rect 16394 12486 16406 12538
rect 16406 12486 16436 12538
rect 16460 12486 16470 12538
rect 16470 12486 16516 12538
rect 16220 12484 16276 12486
rect 16300 12484 16356 12486
rect 16380 12484 16436 12486
rect 16460 12484 16516 12486
rect 13220 10906 13276 10908
rect 13300 10906 13356 10908
rect 13380 10906 13436 10908
rect 13460 10906 13516 10908
rect 13220 10854 13266 10906
rect 13266 10854 13276 10906
rect 13300 10854 13330 10906
rect 13330 10854 13342 10906
rect 13342 10854 13356 10906
rect 13380 10854 13394 10906
rect 13394 10854 13406 10906
rect 13406 10854 13436 10906
rect 13460 10854 13470 10906
rect 13470 10854 13516 10906
rect 13220 10852 13276 10854
rect 13300 10852 13356 10854
rect 13380 10852 13436 10854
rect 13460 10852 13516 10854
rect 16220 11450 16276 11452
rect 16300 11450 16356 11452
rect 16380 11450 16436 11452
rect 16460 11450 16516 11452
rect 16220 11398 16266 11450
rect 16266 11398 16276 11450
rect 16300 11398 16330 11450
rect 16330 11398 16342 11450
rect 16342 11398 16356 11450
rect 16380 11398 16394 11450
rect 16394 11398 16406 11450
rect 16406 11398 16436 11450
rect 16460 11398 16470 11450
rect 16470 11398 16516 11450
rect 16220 11396 16276 11398
rect 16300 11396 16356 11398
rect 16380 11396 16436 11398
rect 16460 11396 16516 11398
rect 13220 9818 13276 9820
rect 13300 9818 13356 9820
rect 13380 9818 13436 9820
rect 13460 9818 13516 9820
rect 13220 9766 13266 9818
rect 13266 9766 13276 9818
rect 13300 9766 13330 9818
rect 13330 9766 13342 9818
rect 13342 9766 13356 9818
rect 13380 9766 13394 9818
rect 13394 9766 13406 9818
rect 13406 9766 13436 9818
rect 13460 9766 13470 9818
rect 13470 9766 13516 9818
rect 13220 9764 13276 9766
rect 13300 9764 13356 9766
rect 13380 9764 13436 9766
rect 13460 9764 13516 9766
rect 16220 10362 16276 10364
rect 16300 10362 16356 10364
rect 16380 10362 16436 10364
rect 16460 10362 16516 10364
rect 16220 10310 16266 10362
rect 16266 10310 16276 10362
rect 16300 10310 16330 10362
rect 16330 10310 16342 10362
rect 16342 10310 16356 10362
rect 16380 10310 16394 10362
rect 16394 10310 16406 10362
rect 16406 10310 16436 10362
rect 16460 10310 16470 10362
rect 16470 10310 16516 10362
rect 16220 10308 16276 10310
rect 16300 10308 16356 10310
rect 16380 10308 16436 10310
rect 16460 10308 16516 10310
rect 19220 20698 19276 20700
rect 19300 20698 19356 20700
rect 19380 20698 19436 20700
rect 19460 20698 19516 20700
rect 19220 20646 19266 20698
rect 19266 20646 19276 20698
rect 19300 20646 19330 20698
rect 19330 20646 19342 20698
rect 19342 20646 19356 20698
rect 19380 20646 19394 20698
rect 19394 20646 19406 20698
rect 19406 20646 19436 20698
rect 19460 20646 19470 20698
rect 19470 20646 19516 20698
rect 19220 20644 19276 20646
rect 19300 20644 19356 20646
rect 19380 20644 19436 20646
rect 19460 20644 19516 20646
rect 19220 19610 19276 19612
rect 19300 19610 19356 19612
rect 19380 19610 19436 19612
rect 19460 19610 19516 19612
rect 19220 19558 19266 19610
rect 19266 19558 19276 19610
rect 19300 19558 19330 19610
rect 19330 19558 19342 19610
rect 19342 19558 19356 19610
rect 19380 19558 19394 19610
rect 19394 19558 19406 19610
rect 19406 19558 19436 19610
rect 19460 19558 19470 19610
rect 19470 19558 19516 19610
rect 19220 19556 19276 19558
rect 19300 19556 19356 19558
rect 19380 19556 19436 19558
rect 19460 19556 19516 19558
rect 19220 18522 19276 18524
rect 19300 18522 19356 18524
rect 19380 18522 19436 18524
rect 19460 18522 19516 18524
rect 19220 18470 19266 18522
rect 19266 18470 19276 18522
rect 19300 18470 19330 18522
rect 19330 18470 19342 18522
rect 19342 18470 19356 18522
rect 19380 18470 19394 18522
rect 19394 18470 19406 18522
rect 19406 18470 19436 18522
rect 19460 18470 19470 18522
rect 19470 18470 19516 18522
rect 19220 18468 19276 18470
rect 19300 18468 19356 18470
rect 19380 18468 19436 18470
rect 19460 18468 19516 18470
rect 19220 17434 19276 17436
rect 19300 17434 19356 17436
rect 19380 17434 19436 17436
rect 19460 17434 19516 17436
rect 19220 17382 19266 17434
rect 19266 17382 19276 17434
rect 19300 17382 19330 17434
rect 19330 17382 19342 17434
rect 19342 17382 19356 17434
rect 19380 17382 19394 17434
rect 19394 17382 19406 17434
rect 19406 17382 19436 17434
rect 19460 17382 19470 17434
rect 19470 17382 19516 17434
rect 19220 17380 19276 17382
rect 19300 17380 19356 17382
rect 19380 17380 19436 17382
rect 19460 17380 19516 17382
rect 20442 21120 20498 21176
rect 19220 16346 19276 16348
rect 19300 16346 19356 16348
rect 19380 16346 19436 16348
rect 19460 16346 19516 16348
rect 19220 16294 19266 16346
rect 19266 16294 19276 16346
rect 19300 16294 19330 16346
rect 19330 16294 19342 16346
rect 19342 16294 19356 16346
rect 19380 16294 19394 16346
rect 19394 16294 19406 16346
rect 19406 16294 19436 16346
rect 19460 16294 19470 16346
rect 19470 16294 19516 16346
rect 19220 16292 19276 16294
rect 19300 16292 19356 16294
rect 19380 16292 19436 16294
rect 19460 16292 19516 16294
rect 19220 15258 19276 15260
rect 19300 15258 19356 15260
rect 19380 15258 19436 15260
rect 19460 15258 19516 15260
rect 19220 15206 19266 15258
rect 19266 15206 19276 15258
rect 19300 15206 19330 15258
rect 19330 15206 19342 15258
rect 19342 15206 19356 15258
rect 19380 15206 19394 15258
rect 19394 15206 19406 15258
rect 19406 15206 19436 15258
rect 19460 15206 19470 15258
rect 19470 15206 19516 15258
rect 19220 15204 19276 15206
rect 19300 15204 19356 15206
rect 19380 15204 19436 15206
rect 19460 15204 19516 15206
rect 19220 14170 19276 14172
rect 19300 14170 19356 14172
rect 19380 14170 19436 14172
rect 19460 14170 19516 14172
rect 19220 14118 19266 14170
rect 19266 14118 19276 14170
rect 19300 14118 19330 14170
rect 19330 14118 19342 14170
rect 19342 14118 19356 14170
rect 19380 14118 19394 14170
rect 19394 14118 19406 14170
rect 19406 14118 19436 14170
rect 19460 14118 19470 14170
rect 19470 14118 19516 14170
rect 19220 14116 19276 14118
rect 19300 14116 19356 14118
rect 19380 14116 19436 14118
rect 19460 14116 19516 14118
rect 20442 15700 20498 15736
rect 20442 15680 20444 15700
rect 20444 15680 20496 15700
rect 20496 15680 20498 15700
rect 19220 13082 19276 13084
rect 19300 13082 19356 13084
rect 19380 13082 19436 13084
rect 19460 13082 19516 13084
rect 19220 13030 19266 13082
rect 19266 13030 19276 13082
rect 19300 13030 19330 13082
rect 19330 13030 19342 13082
rect 19342 13030 19356 13082
rect 19380 13030 19394 13082
rect 19394 13030 19406 13082
rect 19406 13030 19436 13082
rect 19460 13030 19470 13082
rect 19470 13030 19516 13082
rect 19220 13028 19276 13030
rect 19300 13028 19356 13030
rect 19380 13028 19436 13030
rect 19460 13028 19516 13030
rect 19220 11994 19276 11996
rect 19300 11994 19356 11996
rect 19380 11994 19436 11996
rect 19460 11994 19516 11996
rect 19220 11942 19266 11994
rect 19266 11942 19276 11994
rect 19300 11942 19330 11994
rect 19330 11942 19342 11994
rect 19342 11942 19356 11994
rect 19380 11942 19394 11994
rect 19394 11942 19406 11994
rect 19406 11942 19436 11994
rect 19460 11942 19470 11994
rect 19470 11942 19516 11994
rect 19220 11940 19276 11942
rect 19300 11940 19356 11942
rect 19380 11940 19436 11942
rect 19460 11940 19516 11942
rect 10220 8186 10276 8188
rect 10300 8186 10356 8188
rect 10380 8186 10436 8188
rect 10460 8186 10516 8188
rect 10220 8134 10266 8186
rect 10266 8134 10276 8186
rect 10300 8134 10330 8186
rect 10330 8134 10342 8186
rect 10342 8134 10356 8186
rect 10380 8134 10394 8186
rect 10394 8134 10406 8186
rect 10406 8134 10436 8186
rect 10460 8134 10470 8186
rect 10470 8134 10516 8186
rect 10220 8132 10276 8134
rect 10300 8132 10356 8134
rect 10380 8132 10436 8134
rect 10460 8132 10516 8134
rect 13220 8730 13276 8732
rect 13300 8730 13356 8732
rect 13380 8730 13436 8732
rect 13460 8730 13516 8732
rect 13220 8678 13266 8730
rect 13266 8678 13276 8730
rect 13300 8678 13330 8730
rect 13330 8678 13342 8730
rect 13342 8678 13356 8730
rect 13380 8678 13394 8730
rect 13394 8678 13406 8730
rect 13406 8678 13436 8730
rect 13460 8678 13470 8730
rect 13470 8678 13516 8730
rect 13220 8676 13276 8678
rect 13300 8676 13356 8678
rect 13380 8676 13436 8678
rect 13460 8676 13516 8678
rect 10220 7098 10276 7100
rect 10300 7098 10356 7100
rect 10380 7098 10436 7100
rect 10460 7098 10516 7100
rect 10220 7046 10266 7098
rect 10266 7046 10276 7098
rect 10300 7046 10330 7098
rect 10330 7046 10342 7098
rect 10342 7046 10356 7098
rect 10380 7046 10394 7098
rect 10394 7046 10406 7098
rect 10406 7046 10436 7098
rect 10460 7046 10470 7098
rect 10470 7046 10516 7098
rect 10220 7044 10276 7046
rect 10300 7044 10356 7046
rect 10380 7044 10436 7046
rect 10460 7044 10516 7046
rect 10220 6010 10276 6012
rect 10300 6010 10356 6012
rect 10380 6010 10436 6012
rect 10460 6010 10516 6012
rect 10220 5958 10266 6010
rect 10266 5958 10276 6010
rect 10300 5958 10330 6010
rect 10330 5958 10342 6010
rect 10342 5958 10356 6010
rect 10380 5958 10394 6010
rect 10394 5958 10406 6010
rect 10406 5958 10436 6010
rect 10460 5958 10470 6010
rect 10470 5958 10516 6010
rect 10220 5956 10276 5958
rect 10300 5956 10356 5958
rect 10380 5956 10436 5958
rect 10460 5956 10516 5958
rect 10220 4922 10276 4924
rect 10300 4922 10356 4924
rect 10380 4922 10436 4924
rect 10460 4922 10516 4924
rect 10220 4870 10266 4922
rect 10266 4870 10276 4922
rect 10300 4870 10330 4922
rect 10330 4870 10342 4922
rect 10342 4870 10356 4922
rect 10380 4870 10394 4922
rect 10394 4870 10406 4922
rect 10406 4870 10436 4922
rect 10460 4870 10470 4922
rect 10470 4870 10516 4922
rect 10220 4868 10276 4870
rect 10300 4868 10356 4870
rect 10380 4868 10436 4870
rect 10460 4868 10516 4870
rect 9678 3984 9734 4040
rect 10220 3834 10276 3836
rect 10300 3834 10356 3836
rect 10380 3834 10436 3836
rect 10460 3834 10516 3836
rect 10220 3782 10266 3834
rect 10266 3782 10276 3834
rect 10300 3782 10330 3834
rect 10330 3782 10342 3834
rect 10342 3782 10356 3834
rect 10380 3782 10394 3834
rect 10394 3782 10406 3834
rect 10406 3782 10436 3834
rect 10460 3782 10470 3834
rect 10470 3782 10516 3834
rect 10220 3780 10276 3782
rect 10300 3780 10356 3782
rect 10380 3780 10436 3782
rect 10460 3780 10516 3782
rect 13220 7642 13276 7644
rect 13300 7642 13356 7644
rect 13380 7642 13436 7644
rect 13460 7642 13516 7644
rect 13220 7590 13266 7642
rect 13266 7590 13276 7642
rect 13300 7590 13330 7642
rect 13330 7590 13342 7642
rect 13342 7590 13356 7642
rect 13380 7590 13394 7642
rect 13394 7590 13406 7642
rect 13406 7590 13436 7642
rect 13460 7590 13470 7642
rect 13470 7590 13516 7642
rect 13220 7588 13276 7590
rect 13300 7588 13356 7590
rect 13380 7588 13436 7590
rect 13460 7588 13516 7590
rect 13220 6554 13276 6556
rect 13300 6554 13356 6556
rect 13380 6554 13436 6556
rect 13460 6554 13516 6556
rect 13220 6502 13266 6554
rect 13266 6502 13276 6554
rect 13300 6502 13330 6554
rect 13330 6502 13342 6554
rect 13342 6502 13356 6554
rect 13380 6502 13394 6554
rect 13394 6502 13406 6554
rect 13406 6502 13436 6554
rect 13460 6502 13470 6554
rect 13470 6502 13516 6554
rect 13220 6500 13276 6502
rect 13300 6500 13356 6502
rect 13380 6500 13436 6502
rect 13460 6500 13516 6502
rect 13220 5466 13276 5468
rect 13300 5466 13356 5468
rect 13380 5466 13436 5468
rect 13460 5466 13516 5468
rect 13220 5414 13266 5466
rect 13266 5414 13276 5466
rect 13300 5414 13330 5466
rect 13330 5414 13342 5466
rect 13342 5414 13356 5466
rect 13380 5414 13394 5466
rect 13394 5414 13406 5466
rect 13406 5414 13436 5466
rect 13460 5414 13470 5466
rect 13470 5414 13516 5466
rect 13220 5412 13276 5414
rect 13300 5412 13356 5414
rect 13380 5412 13436 5414
rect 13460 5412 13516 5414
rect 16220 9274 16276 9276
rect 16300 9274 16356 9276
rect 16380 9274 16436 9276
rect 16460 9274 16516 9276
rect 16220 9222 16266 9274
rect 16266 9222 16276 9274
rect 16300 9222 16330 9274
rect 16330 9222 16342 9274
rect 16342 9222 16356 9274
rect 16380 9222 16394 9274
rect 16394 9222 16406 9274
rect 16406 9222 16436 9274
rect 16460 9222 16470 9274
rect 16470 9222 16516 9274
rect 16220 9220 16276 9222
rect 16300 9220 16356 9222
rect 16380 9220 16436 9222
rect 16460 9220 16516 9222
rect 16220 8186 16276 8188
rect 16300 8186 16356 8188
rect 16380 8186 16436 8188
rect 16460 8186 16516 8188
rect 16220 8134 16266 8186
rect 16266 8134 16276 8186
rect 16300 8134 16330 8186
rect 16330 8134 16342 8186
rect 16342 8134 16356 8186
rect 16380 8134 16394 8186
rect 16394 8134 16406 8186
rect 16406 8134 16436 8186
rect 16460 8134 16470 8186
rect 16470 8134 16516 8186
rect 16220 8132 16276 8134
rect 16300 8132 16356 8134
rect 16380 8132 16436 8134
rect 16460 8132 16516 8134
rect 16220 7098 16276 7100
rect 16300 7098 16356 7100
rect 16380 7098 16436 7100
rect 16460 7098 16516 7100
rect 16220 7046 16266 7098
rect 16266 7046 16276 7098
rect 16300 7046 16330 7098
rect 16330 7046 16342 7098
rect 16342 7046 16356 7098
rect 16380 7046 16394 7098
rect 16394 7046 16406 7098
rect 16406 7046 16436 7098
rect 16460 7046 16470 7098
rect 16470 7046 16516 7098
rect 16220 7044 16276 7046
rect 16300 7044 16356 7046
rect 16380 7044 16436 7046
rect 16460 7044 16516 7046
rect 16220 6010 16276 6012
rect 16300 6010 16356 6012
rect 16380 6010 16436 6012
rect 16460 6010 16516 6012
rect 16220 5958 16266 6010
rect 16266 5958 16276 6010
rect 16300 5958 16330 6010
rect 16330 5958 16342 6010
rect 16342 5958 16356 6010
rect 16380 5958 16394 6010
rect 16394 5958 16406 6010
rect 16406 5958 16436 6010
rect 16460 5958 16470 6010
rect 16470 5958 16516 6010
rect 16220 5956 16276 5958
rect 16300 5956 16356 5958
rect 16380 5956 16436 5958
rect 16460 5956 16516 5958
rect 19220 10906 19276 10908
rect 19300 10906 19356 10908
rect 19380 10906 19436 10908
rect 19460 10906 19516 10908
rect 19220 10854 19266 10906
rect 19266 10854 19276 10906
rect 19300 10854 19330 10906
rect 19330 10854 19342 10906
rect 19342 10854 19356 10906
rect 19380 10854 19394 10906
rect 19394 10854 19406 10906
rect 19406 10854 19436 10906
rect 19460 10854 19470 10906
rect 19470 10854 19516 10906
rect 19220 10852 19276 10854
rect 19300 10852 19356 10854
rect 19380 10852 19436 10854
rect 19460 10852 19516 10854
rect 19220 9818 19276 9820
rect 19300 9818 19356 9820
rect 19380 9818 19436 9820
rect 19460 9818 19516 9820
rect 19220 9766 19266 9818
rect 19266 9766 19276 9818
rect 19300 9766 19330 9818
rect 19330 9766 19342 9818
rect 19342 9766 19356 9818
rect 19380 9766 19394 9818
rect 19394 9766 19406 9818
rect 19406 9766 19436 9818
rect 19460 9766 19470 9818
rect 19470 9766 19516 9818
rect 19220 9764 19276 9766
rect 19300 9764 19356 9766
rect 19380 9764 19436 9766
rect 19460 9764 19516 9766
rect 20442 10240 20498 10296
rect 19220 8730 19276 8732
rect 19300 8730 19356 8732
rect 19380 8730 19436 8732
rect 19460 8730 19516 8732
rect 19220 8678 19266 8730
rect 19266 8678 19276 8730
rect 19300 8678 19330 8730
rect 19330 8678 19342 8730
rect 19342 8678 19356 8730
rect 19380 8678 19394 8730
rect 19394 8678 19406 8730
rect 19406 8678 19436 8730
rect 19460 8678 19470 8730
rect 19470 8678 19516 8730
rect 19220 8676 19276 8678
rect 19300 8676 19356 8678
rect 19380 8676 19436 8678
rect 19460 8676 19516 8678
rect 19220 7642 19276 7644
rect 19300 7642 19356 7644
rect 19380 7642 19436 7644
rect 19460 7642 19516 7644
rect 19220 7590 19266 7642
rect 19266 7590 19276 7642
rect 19300 7590 19330 7642
rect 19330 7590 19342 7642
rect 19342 7590 19356 7642
rect 19380 7590 19394 7642
rect 19394 7590 19406 7642
rect 19406 7590 19436 7642
rect 19460 7590 19470 7642
rect 19470 7590 19516 7642
rect 19220 7588 19276 7590
rect 19300 7588 19356 7590
rect 19380 7588 19436 7590
rect 19460 7588 19516 7590
rect 19220 6554 19276 6556
rect 19300 6554 19356 6556
rect 19380 6554 19436 6556
rect 19460 6554 19516 6556
rect 19220 6502 19266 6554
rect 19266 6502 19276 6554
rect 19300 6502 19330 6554
rect 19330 6502 19342 6554
rect 19342 6502 19356 6554
rect 19380 6502 19394 6554
rect 19394 6502 19406 6554
rect 19406 6502 19436 6554
rect 19460 6502 19470 6554
rect 19470 6502 19516 6554
rect 19220 6500 19276 6502
rect 19300 6500 19356 6502
rect 19380 6500 19436 6502
rect 19460 6500 19516 6502
rect 19220 5466 19276 5468
rect 19300 5466 19356 5468
rect 19380 5466 19436 5468
rect 19460 5466 19516 5468
rect 19220 5414 19266 5466
rect 19266 5414 19276 5466
rect 19300 5414 19330 5466
rect 19330 5414 19342 5466
rect 19342 5414 19356 5466
rect 19380 5414 19394 5466
rect 19394 5414 19406 5466
rect 19406 5414 19436 5466
rect 19460 5414 19470 5466
rect 19470 5414 19516 5466
rect 19220 5412 19276 5414
rect 19300 5412 19356 5414
rect 19380 5412 19436 5414
rect 19460 5412 19516 5414
rect 16220 4922 16276 4924
rect 16300 4922 16356 4924
rect 16380 4922 16436 4924
rect 16460 4922 16516 4924
rect 16220 4870 16266 4922
rect 16266 4870 16276 4922
rect 16300 4870 16330 4922
rect 16330 4870 16342 4922
rect 16342 4870 16356 4922
rect 16380 4870 16394 4922
rect 16394 4870 16406 4922
rect 16406 4870 16436 4922
rect 16460 4870 16470 4922
rect 16470 4870 16516 4922
rect 16220 4868 16276 4870
rect 16300 4868 16356 4870
rect 16380 4868 16436 4870
rect 16460 4868 16516 4870
rect 13220 4378 13276 4380
rect 13300 4378 13356 4380
rect 13380 4378 13436 4380
rect 13460 4378 13516 4380
rect 13220 4326 13266 4378
rect 13266 4326 13276 4378
rect 13300 4326 13330 4378
rect 13330 4326 13342 4378
rect 13342 4326 13356 4378
rect 13380 4326 13394 4378
rect 13394 4326 13406 4378
rect 13406 4326 13436 4378
rect 13460 4326 13470 4378
rect 13470 4326 13516 4378
rect 13220 4324 13276 4326
rect 13300 4324 13356 4326
rect 13380 4324 13436 4326
rect 13460 4324 13516 4326
rect 10220 2746 10276 2748
rect 10300 2746 10356 2748
rect 10380 2746 10436 2748
rect 10460 2746 10516 2748
rect 10220 2694 10266 2746
rect 10266 2694 10276 2746
rect 10300 2694 10330 2746
rect 10330 2694 10342 2746
rect 10342 2694 10356 2746
rect 10380 2694 10394 2746
rect 10394 2694 10406 2746
rect 10406 2694 10436 2746
rect 10460 2694 10470 2746
rect 10470 2694 10516 2746
rect 10220 2692 10276 2694
rect 10300 2692 10356 2694
rect 10380 2692 10436 2694
rect 10460 2692 10516 2694
rect 13220 3290 13276 3292
rect 13300 3290 13356 3292
rect 13380 3290 13436 3292
rect 13460 3290 13516 3292
rect 13220 3238 13266 3290
rect 13266 3238 13276 3290
rect 13300 3238 13330 3290
rect 13330 3238 13342 3290
rect 13342 3238 13356 3290
rect 13380 3238 13394 3290
rect 13394 3238 13406 3290
rect 13406 3238 13436 3290
rect 13460 3238 13470 3290
rect 13470 3238 13516 3290
rect 13220 3236 13276 3238
rect 13300 3236 13356 3238
rect 13380 3236 13436 3238
rect 13460 3236 13516 3238
rect 20810 4800 20866 4856
rect 19220 4378 19276 4380
rect 19300 4378 19356 4380
rect 19380 4378 19436 4380
rect 19460 4378 19516 4380
rect 19220 4326 19266 4378
rect 19266 4326 19276 4378
rect 19300 4326 19330 4378
rect 19330 4326 19342 4378
rect 19342 4326 19356 4378
rect 19380 4326 19394 4378
rect 19394 4326 19406 4378
rect 19406 4326 19436 4378
rect 19460 4326 19470 4378
rect 19470 4326 19516 4378
rect 19220 4324 19276 4326
rect 19300 4324 19356 4326
rect 19380 4324 19436 4326
rect 19460 4324 19516 4326
rect 16220 3834 16276 3836
rect 16300 3834 16356 3836
rect 16380 3834 16436 3836
rect 16460 3834 16516 3836
rect 16220 3782 16266 3834
rect 16266 3782 16276 3834
rect 16300 3782 16330 3834
rect 16330 3782 16342 3834
rect 16342 3782 16356 3834
rect 16380 3782 16394 3834
rect 16394 3782 16406 3834
rect 16406 3782 16436 3834
rect 16460 3782 16470 3834
rect 16470 3782 16516 3834
rect 16220 3780 16276 3782
rect 16300 3780 16356 3782
rect 16380 3780 16436 3782
rect 16460 3780 16516 3782
rect 19220 3290 19276 3292
rect 19300 3290 19356 3292
rect 19380 3290 19436 3292
rect 19460 3290 19516 3292
rect 19220 3238 19266 3290
rect 19266 3238 19276 3290
rect 19300 3238 19330 3290
rect 19330 3238 19342 3290
rect 19342 3238 19356 3290
rect 19380 3238 19394 3290
rect 19394 3238 19406 3290
rect 19406 3238 19436 3290
rect 19460 3238 19470 3290
rect 19470 3238 19516 3290
rect 19220 3236 19276 3238
rect 19300 3236 19356 3238
rect 19380 3236 19436 3238
rect 19460 3236 19516 3238
rect 16220 2746 16276 2748
rect 16300 2746 16356 2748
rect 16380 2746 16436 2748
rect 16460 2746 16516 2748
rect 16220 2694 16266 2746
rect 16266 2694 16276 2746
rect 16300 2694 16330 2746
rect 16330 2694 16342 2746
rect 16342 2694 16356 2746
rect 16380 2694 16394 2746
rect 16394 2694 16406 2746
rect 16406 2694 16436 2746
rect 16460 2694 16470 2746
rect 16470 2694 16516 2746
rect 16220 2692 16276 2694
rect 16300 2692 16356 2694
rect 16380 2692 16436 2694
rect 16460 2692 16516 2694
rect 7220 2202 7276 2204
rect 7300 2202 7356 2204
rect 7380 2202 7436 2204
rect 7460 2202 7516 2204
rect 7220 2150 7266 2202
rect 7266 2150 7276 2202
rect 7300 2150 7330 2202
rect 7330 2150 7342 2202
rect 7342 2150 7356 2202
rect 7380 2150 7394 2202
rect 7394 2150 7406 2202
rect 7406 2150 7436 2202
rect 7460 2150 7470 2202
rect 7470 2150 7516 2202
rect 7220 2148 7276 2150
rect 7300 2148 7356 2150
rect 7380 2148 7436 2150
rect 7460 2148 7516 2150
rect 13220 2202 13276 2204
rect 13300 2202 13356 2204
rect 13380 2202 13436 2204
rect 13460 2202 13516 2204
rect 13220 2150 13266 2202
rect 13266 2150 13276 2202
rect 13300 2150 13330 2202
rect 13330 2150 13342 2202
rect 13342 2150 13356 2202
rect 13380 2150 13394 2202
rect 13394 2150 13406 2202
rect 13406 2150 13436 2202
rect 13460 2150 13470 2202
rect 13470 2150 13516 2202
rect 13220 2148 13276 2150
rect 13300 2148 13356 2150
rect 13380 2148 13436 2150
rect 13460 2148 13516 2150
rect 19220 2202 19276 2204
rect 19300 2202 19356 2204
rect 19380 2202 19436 2204
rect 19460 2202 19516 2204
rect 19220 2150 19266 2202
rect 19266 2150 19276 2202
rect 19300 2150 19330 2202
rect 19330 2150 19342 2202
rect 19342 2150 19356 2202
rect 19380 2150 19394 2202
rect 19394 2150 19406 2202
rect 19406 2150 19436 2202
rect 19460 2150 19470 2202
rect 19470 2150 19516 2202
rect 19220 2148 19276 2150
rect 19300 2148 19356 2150
rect 19380 2148 19436 2150
rect 19460 2148 19516 2150
<< metal3 >>
rect 0 21858 800 21888
rect 3141 21858 3207 21861
rect 0 21856 3207 21858
rect 0 21800 3146 21856
rect 3202 21800 3207 21856
rect 0 21798 3207 21800
rect 0 21768 800 21798
rect 3141 21795 3207 21798
rect 7210 21792 7526 21793
rect 7210 21728 7216 21792
rect 7280 21728 7296 21792
rect 7360 21728 7376 21792
rect 7440 21728 7456 21792
rect 7520 21728 7526 21792
rect 7210 21727 7526 21728
rect 13210 21792 13526 21793
rect 13210 21728 13216 21792
rect 13280 21728 13296 21792
rect 13360 21728 13376 21792
rect 13440 21728 13456 21792
rect 13520 21728 13526 21792
rect 13210 21727 13526 21728
rect 19210 21792 19526 21793
rect 19210 21728 19216 21792
rect 19280 21728 19296 21792
rect 19360 21728 19376 21792
rect 19440 21728 19456 21792
rect 19520 21728 19526 21792
rect 19210 21727 19526 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 10210 21248 10526 21249
rect 10210 21184 10216 21248
rect 10280 21184 10296 21248
rect 10360 21184 10376 21248
rect 10440 21184 10456 21248
rect 10520 21184 10526 21248
rect 10210 21183 10526 21184
rect 16210 21248 16526 21249
rect 16210 21184 16216 21248
rect 16280 21184 16296 21248
rect 16360 21184 16376 21248
rect 16440 21184 16456 21248
rect 16520 21184 16526 21248
rect 16210 21183 16526 21184
rect 20437 21178 20503 21181
rect 21118 21178 21918 21208
rect 20437 21176 21918 21178
rect 20437 21120 20442 21176
rect 20498 21120 21918 21176
rect 20437 21118 21918 21120
rect 20437 21115 20503 21118
rect 21118 21088 21918 21118
rect 7210 20704 7526 20705
rect 7210 20640 7216 20704
rect 7280 20640 7296 20704
rect 7360 20640 7376 20704
rect 7440 20640 7456 20704
rect 7520 20640 7526 20704
rect 7210 20639 7526 20640
rect 13210 20704 13526 20705
rect 13210 20640 13216 20704
rect 13280 20640 13296 20704
rect 13360 20640 13376 20704
rect 13440 20640 13456 20704
rect 13520 20640 13526 20704
rect 13210 20639 13526 20640
rect 19210 20704 19526 20705
rect 19210 20640 19216 20704
rect 19280 20640 19296 20704
rect 19360 20640 19376 20704
rect 19440 20640 19456 20704
rect 19520 20640 19526 20704
rect 19210 20639 19526 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 10210 20160 10526 20161
rect 10210 20096 10216 20160
rect 10280 20096 10296 20160
rect 10360 20096 10376 20160
rect 10440 20096 10456 20160
rect 10520 20096 10526 20160
rect 10210 20095 10526 20096
rect 16210 20160 16526 20161
rect 16210 20096 16216 20160
rect 16280 20096 16296 20160
rect 16360 20096 16376 20160
rect 16440 20096 16456 20160
rect 16520 20096 16526 20160
rect 16210 20095 16526 20096
rect 7210 19616 7526 19617
rect 7210 19552 7216 19616
rect 7280 19552 7296 19616
rect 7360 19552 7376 19616
rect 7440 19552 7456 19616
rect 7520 19552 7526 19616
rect 7210 19551 7526 19552
rect 13210 19616 13526 19617
rect 13210 19552 13216 19616
rect 13280 19552 13296 19616
rect 13360 19552 13376 19616
rect 13440 19552 13456 19616
rect 13520 19552 13526 19616
rect 13210 19551 13526 19552
rect 19210 19616 19526 19617
rect 19210 19552 19216 19616
rect 19280 19552 19296 19616
rect 19360 19552 19376 19616
rect 19440 19552 19456 19616
rect 19520 19552 19526 19616
rect 19210 19551 19526 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 10210 19072 10526 19073
rect 10210 19008 10216 19072
rect 10280 19008 10296 19072
rect 10360 19008 10376 19072
rect 10440 19008 10456 19072
rect 10520 19008 10526 19072
rect 10210 19007 10526 19008
rect 16210 19072 16526 19073
rect 16210 19008 16216 19072
rect 16280 19008 16296 19072
rect 16360 19008 16376 19072
rect 16440 19008 16456 19072
rect 16520 19008 16526 19072
rect 16210 19007 16526 19008
rect 7210 18528 7526 18529
rect 7210 18464 7216 18528
rect 7280 18464 7296 18528
rect 7360 18464 7376 18528
rect 7440 18464 7456 18528
rect 7520 18464 7526 18528
rect 7210 18463 7526 18464
rect 13210 18528 13526 18529
rect 13210 18464 13216 18528
rect 13280 18464 13296 18528
rect 13360 18464 13376 18528
rect 13440 18464 13456 18528
rect 13520 18464 13526 18528
rect 13210 18463 13526 18464
rect 19210 18528 19526 18529
rect 19210 18464 19216 18528
rect 19280 18464 19296 18528
rect 19360 18464 19376 18528
rect 19440 18464 19456 18528
rect 19520 18464 19526 18528
rect 19210 18463 19526 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 10210 17984 10526 17985
rect 10210 17920 10216 17984
rect 10280 17920 10296 17984
rect 10360 17920 10376 17984
rect 10440 17920 10456 17984
rect 10520 17920 10526 17984
rect 10210 17919 10526 17920
rect 16210 17984 16526 17985
rect 16210 17920 16216 17984
rect 16280 17920 16296 17984
rect 16360 17920 16376 17984
rect 16440 17920 16456 17984
rect 16520 17920 16526 17984
rect 16210 17919 16526 17920
rect 7210 17440 7526 17441
rect 7210 17376 7216 17440
rect 7280 17376 7296 17440
rect 7360 17376 7376 17440
rect 7440 17376 7456 17440
rect 7520 17376 7526 17440
rect 7210 17375 7526 17376
rect 13210 17440 13526 17441
rect 13210 17376 13216 17440
rect 13280 17376 13296 17440
rect 13360 17376 13376 17440
rect 13440 17376 13456 17440
rect 13520 17376 13526 17440
rect 13210 17375 13526 17376
rect 19210 17440 19526 17441
rect 19210 17376 19216 17440
rect 19280 17376 19296 17440
rect 19360 17376 19376 17440
rect 19440 17376 19456 17440
rect 19520 17376 19526 17440
rect 19210 17375 19526 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 10210 16896 10526 16897
rect 10210 16832 10216 16896
rect 10280 16832 10296 16896
rect 10360 16832 10376 16896
rect 10440 16832 10456 16896
rect 10520 16832 10526 16896
rect 10210 16831 10526 16832
rect 16210 16896 16526 16897
rect 16210 16832 16216 16896
rect 16280 16832 16296 16896
rect 16360 16832 16376 16896
rect 16440 16832 16456 16896
rect 16520 16832 16526 16896
rect 16210 16831 16526 16832
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 7210 16352 7526 16353
rect 7210 16288 7216 16352
rect 7280 16288 7296 16352
rect 7360 16288 7376 16352
rect 7440 16288 7456 16352
rect 7520 16288 7526 16352
rect 7210 16287 7526 16288
rect 13210 16352 13526 16353
rect 13210 16288 13216 16352
rect 13280 16288 13296 16352
rect 13360 16288 13376 16352
rect 13440 16288 13456 16352
rect 13520 16288 13526 16352
rect 13210 16287 13526 16288
rect 19210 16352 19526 16353
rect 19210 16288 19216 16352
rect 19280 16288 19296 16352
rect 19360 16288 19376 16352
rect 19440 16288 19456 16352
rect 19520 16288 19526 16352
rect 19210 16287 19526 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 10210 15808 10526 15809
rect 10210 15744 10216 15808
rect 10280 15744 10296 15808
rect 10360 15744 10376 15808
rect 10440 15744 10456 15808
rect 10520 15744 10526 15808
rect 10210 15743 10526 15744
rect 16210 15808 16526 15809
rect 16210 15744 16216 15808
rect 16280 15744 16296 15808
rect 16360 15744 16376 15808
rect 16440 15744 16456 15808
rect 16520 15744 16526 15808
rect 16210 15743 16526 15744
rect 20437 15738 20503 15741
rect 21118 15738 21918 15768
rect 20437 15736 21918 15738
rect 20437 15680 20442 15736
rect 20498 15680 21918 15736
rect 20437 15678 21918 15680
rect 20437 15675 20503 15678
rect 21118 15648 21918 15678
rect 7210 15264 7526 15265
rect 7210 15200 7216 15264
rect 7280 15200 7296 15264
rect 7360 15200 7376 15264
rect 7440 15200 7456 15264
rect 7520 15200 7526 15264
rect 7210 15199 7526 15200
rect 13210 15264 13526 15265
rect 13210 15200 13216 15264
rect 13280 15200 13296 15264
rect 13360 15200 13376 15264
rect 13440 15200 13456 15264
rect 13520 15200 13526 15264
rect 13210 15199 13526 15200
rect 19210 15264 19526 15265
rect 19210 15200 19216 15264
rect 19280 15200 19296 15264
rect 19360 15200 19376 15264
rect 19440 15200 19456 15264
rect 19520 15200 19526 15264
rect 19210 15199 19526 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 10210 14720 10526 14721
rect 10210 14656 10216 14720
rect 10280 14656 10296 14720
rect 10360 14656 10376 14720
rect 10440 14656 10456 14720
rect 10520 14656 10526 14720
rect 10210 14655 10526 14656
rect 16210 14720 16526 14721
rect 16210 14656 16216 14720
rect 16280 14656 16296 14720
rect 16360 14656 16376 14720
rect 16440 14656 16456 14720
rect 16520 14656 16526 14720
rect 16210 14655 16526 14656
rect 7210 14176 7526 14177
rect 7210 14112 7216 14176
rect 7280 14112 7296 14176
rect 7360 14112 7376 14176
rect 7440 14112 7456 14176
rect 7520 14112 7526 14176
rect 7210 14111 7526 14112
rect 13210 14176 13526 14177
rect 13210 14112 13216 14176
rect 13280 14112 13296 14176
rect 13360 14112 13376 14176
rect 13440 14112 13456 14176
rect 13520 14112 13526 14176
rect 13210 14111 13526 14112
rect 19210 14176 19526 14177
rect 19210 14112 19216 14176
rect 19280 14112 19296 14176
rect 19360 14112 19376 14176
rect 19440 14112 19456 14176
rect 19520 14112 19526 14176
rect 19210 14111 19526 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 10210 13632 10526 13633
rect 10210 13568 10216 13632
rect 10280 13568 10296 13632
rect 10360 13568 10376 13632
rect 10440 13568 10456 13632
rect 10520 13568 10526 13632
rect 10210 13567 10526 13568
rect 16210 13632 16526 13633
rect 16210 13568 16216 13632
rect 16280 13568 16296 13632
rect 16360 13568 16376 13632
rect 16440 13568 16456 13632
rect 16520 13568 16526 13632
rect 16210 13567 16526 13568
rect 7210 13088 7526 13089
rect 7210 13024 7216 13088
rect 7280 13024 7296 13088
rect 7360 13024 7376 13088
rect 7440 13024 7456 13088
rect 7520 13024 7526 13088
rect 7210 13023 7526 13024
rect 13210 13088 13526 13089
rect 13210 13024 13216 13088
rect 13280 13024 13296 13088
rect 13360 13024 13376 13088
rect 13440 13024 13456 13088
rect 13520 13024 13526 13088
rect 13210 13023 13526 13024
rect 19210 13088 19526 13089
rect 19210 13024 19216 13088
rect 19280 13024 19296 13088
rect 19360 13024 19376 13088
rect 19440 13024 19456 13088
rect 19520 13024 19526 13088
rect 19210 13023 19526 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 10210 12544 10526 12545
rect 10210 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10526 12544
rect 10210 12479 10526 12480
rect 16210 12544 16526 12545
rect 16210 12480 16216 12544
rect 16280 12480 16296 12544
rect 16360 12480 16376 12544
rect 16440 12480 16456 12544
rect 16520 12480 16526 12544
rect 16210 12479 16526 12480
rect 7210 12000 7526 12001
rect 7210 11936 7216 12000
rect 7280 11936 7296 12000
rect 7360 11936 7376 12000
rect 7440 11936 7456 12000
rect 7520 11936 7526 12000
rect 7210 11935 7526 11936
rect 13210 12000 13526 12001
rect 13210 11936 13216 12000
rect 13280 11936 13296 12000
rect 13360 11936 13376 12000
rect 13440 11936 13456 12000
rect 13520 11936 13526 12000
rect 13210 11935 13526 11936
rect 19210 12000 19526 12001
rect 19210 11936 19216 12000
rect 19280 11936 19296 12000
rect 19360 11936 19376 12000
rect 19440 11936 19456 12000
rect 19520 11936 19526 12000
rect 19210 11935 19526 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 10210 11456 10526 11457
rect 10210 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10526 11456
rect 10210 11391 10526 11392
rect 16210 11456 16526 11457
rect 16210 11392 16216 11456
rect 16280 11392 16296 11456
rect 16360 11392 16376 11456
rect 16440 11392 16456 11456
rect 16520 11392 16526 11456
rect 16210 11391 16526 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 7210 10912 7526 10913
rect 7210 10848 7216 10912
rect 7280 10848 7296 10912
rect 7360 10848 7376 10912
rect 7440 10848 7456 10912
rect 7520 10848 7526 10912
rect 7210 10847 7526 10848
rect 13210 10912 13526 10913
rect 13210 10848 13216 10912
rect 13280 10848 13296 10912
rect 13360 10848 13376 10912
rect 13440 10848 13456 10912
rect 13520 10848 13526 10912
rect 13210 10847 13526 10848
rect 19210 10912 19526 10913
rect 19210 10848 19216 10912
rect 19280 10848 19296 10912
rect 19360 10848 19376 10912
rect 19440 10848 19456 10912
rect 19520 10848 19526 10912
rect 19210 10847 19526 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 10210 10368 10526 10369
rect 10210 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10526 10368
rect 10210 10303 10526 10304
rect 16210 10368 16526 10369
rect 16210 10304 16216 10368
rect 16280 10304 16296 10368
rect 16360 10304 16376 10368
rect 16440 10304 16456 10368
rect 16520 10304 16526 10368
rect 16210 10303 16526 10304
rect 20437 10298 20503 10301
rect 21118 10298 21918 10328
rect 20437 10296 21918 10298
rect 20437 10240 20442 10296
rect 20498 10240 21918 10296
rect 20437 10238 21918 10240
rect 20437 10235 20503 10238
rect 21118 10208 21918 10238
rect 7210 9824 7526 9825
rect 7210 9760 7216 9824
rect 7280 9760 7296 9824
rect 7360 9760 7376 9824
rect 7440 9760 7456 9824
rect 7520 9760 7526 9824
rect 7210 9759 7526 9760
rect 13210 9824 13526 9825
rect 13210 9760 13216 9824
rect 13280 9760 13296 9824
rect 13360 9760 13376 9824
rect 13440 9760 13456 9824
rect 13520 9760 13526 9824
rect 13210 9759 13526 9760
rect 19210 9824 19526 9825
rect 19210 9760 19216 9824
rect 19280 9760 19296 9824
rect 19360 9760 19376 9824
rect 19440 9760 19456 9824
rect 19520 9760 19526 9824
rect 19210 9759 19526 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 10210 9280 10526 9281
rect 10210 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10526 9280
rect 10210 9215 10526 9216
rect 16210 9280 16526 9281
rect 16210 9216 16216 9280
rect 16280 9216 16296 9280
rect 16360 9216 16376 9280
rect 16440 9216 16456 9280
rect 16520 9216 16526 9280
rect 16210 9215 16526 9216
rect 7210 8736 7526 8737
rect 7210 8672 7216 8736
rect 7280 8672 7296 8736
rect 7360 8672 7376 8736
rect 7440 8672 7456 8736
rect 7520 8672 7526 8736
rect 7210 8671 7526 8672
rect 13210 8736 13526 8737
rect 13210 8672 13216 8736
rect 13280 8672 13296 8736
rect 13360 8672 13376 8736
rect 13440 8672 13456 8736
rect 13520 8672 13526 8736
rect 13210 8671 13526 8672
rect 19210 8736 19526 8737
rect 19210 8672 19216 8736
rect 19280 8672 19296 8736
rect 19360 8672 19376 8736
rect 19440 8672 19456 8736
rect 19520 8672 19526 8736
rect 19210 8671 19526 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 10210 8192 10526 8193
rect 10210 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10526 8192
rect 10210 8127 10526 8128
rect 16210 8192 16526 8193
rect 16210 8128 16216 8192
rect 16280 8128 16296 8192
rect 16360 8128 16376 8192
rect 16440 8128 16456 8192
rect 16520 8128 16526 8192
rect 16210 8127 16526 8128
rect 7210 7648 7526 7649
rect 7210 7584 7216 7648
rect 7280 7584 7296 7648
rect 7360 7584 7376 7648
rect 7440 7584 7456 7648
rect 7520 7584 7526 7648
rect 7210 7583 7526 7584
rect 13210 7648 13526 7649
rect 13210 7584 13216 7648
rect 13280 7584 13296 7648
rect 13360 7584 13376 7648
rect 13440 7584 13456 7648
rect 13520 7584 13526 7648
rect 13210 7583 13526 7584
rect 19210 7648 19526 7649
rect 19210 7584 19216 7648
rect 19280 7584 19296 7648
rect 19360 7584 19376 7648
rect 19440 7584 19456 7648
rect 19520 7584 19526 7648
rect 19210 7583 19526 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 10210 7104 10526 7105
rect 10210 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10526 7104
rect 10210 7039 10526 7040
rect 16210 7104 16526 7105
rect 16210 7040 16216 7104
rect 16280 7040 16296 7104
rect 16360 7040 16376 7104
rect 16440 7040 16456 7104
rect 16520 7040 16526 7104
rect 16210 7039 16526 7040
rect 7210 6560 7526 6561
rect 7210 6496 7216 6560
rect 7280 6496 7296 6560
rect 7360 6496 7376 6560
rect 7440 6496 7456 6560
rect 7520 6496 7526 6560
rect 7210 6495 7526 6496
rect 13210 6560 13526 6561
rect 13210 6496 13216 6560
rect 13280 6496 13296 6560
rect 13360 6496 13376 6560
rect 13440 6496 13456 6560
rect 13520 6496 13526 6560
rect 13210 6495 13526 6496
rect 19210 6560 19526 6561
rect 19210 6496 19216 6560
rect 19280 6496 19296 6560
rect 19360 6496 19376 6560
rect 19440 6496 19456 6560
rect 19520 6496 19526 6560
rect 19210 6495 19526 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 10210 6016 10526 6017
rect 10210 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10526 6016
rect 10210 5951 10526 5952
rect 16210 6016 16526 6017
rect 16210 5952 16216 6016
rect 16280 5952 16296 6016
rect 16360 5952 16376 6016
rect 16440 5952 16456 6016
rect 16520 5952 16526 6016
rect 16210 5951 16526 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 7210 5472 7526 5473
rect 7210 5408 7216 5472
rect 7280 5408 7296 5472
rect 7360 5408 7376 5472
rect 7440 5408 7456 5472
rect 7520 5408 7526 5472
rect 7210 5407 7526 5408
rect 13210 5472 13526 5473
rect 13210 5408 13216 5472
rect 13280 5408 13296 5472
rect 13360 5408 13376 5472
rect 13440 5408 13456 5472
rect 13520 5408 13526 5472
rect 13210 5407 13526 5408
rect 19210 5472 19526 5473
rect 19210 5408 19216 5472
rect 19280 5408 19296 5472
rect 19360 5408 19376 5472
rect 19440 5408 19456 5472
rect 19520 5408 19526 5472
rect 19210 5407 19526 5408
rect 6269 5266 6335 5269
rect 7097 5266 7163 5269
rect 6269 5264 7163 5266
rect 6269 5208 6274 5264
rect 6330 5208 7102 5264
rect 7158 5208 7163 5264
rect 6269 5206 7163 5208
rect 6269 5203 6335 5206
rect 7097 5203 7163 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 10210 4928 10526 4929
rect 10210 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10526 4928
rect 10210 4863 10526 4864
rect 16210 4928 16526 4929
rect 16210 4864 16216 4928
rect 16280 4864 16296 4928
rect 16360 4864 16376 4928
rect 16440 4864 16456 4928
rect 16520 4864 16526 4928
rect 16210 4863 16526 4864
rect 20805 4858 20871 4861
rect 21118 4858 21918 4888
rect 20805 4856 21918 4858
rect 20805 4800 20810 4856
rect 20866 4800 21918 4856
rect 20805 4798 21918 4800
rect 20805 4795 20871 4798
rect 21118 4768 21918 4798
rect 7210 4384 7526 4385
rect 7210 4320 7216 4384
rect 7280 4320 7296 4384
rect 7360 4320 7376 4384
rect 7440 4320 7456 4384
rect 7520 4320 7526 4384
rect 7210 4319 7526 4320
rect 13210 4384 13526 4385
rect 13210 4320 13216 4384
rect 13280 4320 13296 4384
rect 13360 4320 13376 4384
rect 13440 4320 13456 4384
rect 13520 4320 13526 4384
rect 13210 4319 13526 4320
rect 19210 4384 19526 4385
rect 19210 4320 19216 4384
rect 19280 4320 19296 4384
rect 19360 4320 19376 4384
rect 19440 4320 19456 4384
rect 19520 4320 19526 4384
rect 19210 4319 19526 4320
rect 7649 4042 7715 4045
rect 9673 4042 9739 4045
rect 7649 4040 9739 4042
rect 7649 3984 7654 4040
rect 7710 3984 9678 4040
rect 9734 3984 9739 4040
rect 7649 3982 9739 3984
rect 7649 3979 7715 3982
rect 9673 3979 9739 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 10210 3840 10526 3841
rect 10210 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10526 3840
rect 10210 3775 10526 3776
rect 16210 3840 16526 3841
rect 16210 3776 16216 3840
rect 16280 3776 16296 3840
rect 16360 3776 16376 3840
rect 16440 3776 16456 3840
rect 16520 3776 16526 3840
rect 16210 3775 16526 3776
rect 7210 3296 7526 3297
rect 7210 3232 7216 3296
rect 7280 3232 7296 3296
rect 7360 3232 7376 3296
rect 7440 3232 7456 3296
rect 7520 3232 7526 3296
rect 7210 3231 7526 3232
rect 13210 3296 13526 3297
rect 13210 3232 13216 3296
rect 13280 3232 13296 3296
rect 13360 3232 13376 3296
rect 13440 3232 13456 3296
rect 13520 3232 13526 3296
rect 13210 3231 13526 3232
rect 19210 3296 19526 3297
rect 19210 3232 19216 3296
rect 19280 3232 19296 3296
rect 19360 3232 19376 3296
rect 19440 3232 19456 3296
rect 19520 3232 19526 3296
rect 19210 3231 19526 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 10210 2752 10526 2753
rect 10210 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10526 2752
rect 10210 2687 10526 2688
rect 16210 2752 16526 2753
rect 16210 2688 16216 2752
rect 16280 2688 16296 2752
rect 16360 2688 16376 2752
rect 16440 2688 16456 2752
rect 16520 2688 16526 2752
rect 16210 2687 16526 2688
rect 7210 2208 7526 2209
rect 7210 2144 7216 2208
rect 7280 2144 7296 2208
rect 7360 2144 7376 2208
rect 7440 2144 7456 2208
rect 7520 2144 7526 2208
rect 7210 2143 7526 2144
rect 13210 2208 13526 2209
rect 13210 2144 13216 2208
rect 13280 2144 13296 2208
rect 13360 2144 13376 2208
rect 13440 2144 13456 2208
rect 13520 2144 13526 2208
rect 13210 2143 13526 2144
rect 19210 2208 19526 2209
rect 19210 2144 19216 2208
rect 19280 2144 19296 2208
rect 19360 2144 19376 2208
rect 19440 2144 19456 2208
rect 19520 2144 19526 2208
rect 19210 2143 19526 2144
<< via3 >>
rect 7216 21788 7280 21792
rect 7216 21732 7220 21788
rect 7220 21732 7276 21788
rect 7276 21732 7280 21788
rect 7216 21728 7280 21732
rect 7296 21788 7360 21792
rect 7296 21732 7300 21788
rect 7300 21732 7356 21788
rect 7356 21732 7360 21788
rect 7296 21728 7360 21732
rect 7376 21788 7440 21792
rect 7376 21732 7380 21788
rect 7380 21732 7436 21788
rect 7436 21732 7440 21788
rect 7376 21728 7440 21732
rect 7456 21788 7520 21792
rect 7456 21732 7460 21788
rect 7460 21732 7516 21788
rect 7516 21732 7520 21788
rect 7456 21728 7520 21732
rect 13216 21788 13280 21792
rect 13216 21732 13220 21788
rect 13220 21732 13276 21788
rect 13276 21732 13280 21788
rect 13216 21728 13280 21732
rect 13296 21788 13360 21792
rect 13296 21732 13300 21788
rect 13300 21732 13356 21788
rect 13356 21732 13360 21788
rect 13296 21728 13360 21732
rect 13376 21788 13440 21792
rect 13376 21732 13380 21788
rect 13380 21732 13436 21788
rect 13436 21732 13440 21788
rect 13376 21728 13440 21732
rect 13456 21788 13520 21792
rect 13456 21732 13460 21788
rect 13460 21732 13516 21788
rect 13516 21732 13520 21788
rect 13456 21728 13520 21732
rect 19216 21788 19280 21792
rect 19216 21732 19220 21788
rect 19220 21732 19276 21788
rect 19276 21732 19280 21788
rect 19216 21728 19280 21732
rect 19296 21788 19360 21792
rect 19296 21732 19300 21788
rect 19300 21732 19356 21788
rect 19356 21732 19360 21788
rect 19296 21728 19360 21732
rect 19376 21788 19440 21792
rect 19376 21732 19380 21788
rect 19380 21732 19436 21788
rect 19436 21732 19440 21788
rect 19376 21728 19440 21732
rect 19456 21788 19520 21792
rect 19456 21732 19460 21788
rect 19460 21732 19516 21788
rect 19516 21732 19520 21788
rect 19456 21728 19520 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 10216 21244 10280 21248
rect 10216 21188 10220 21244
rect 10220 21188 10276 21244
rect 10276 21188 10280 21244
rect 10216 21184 10280 21188
rect 10296 21244 10360 21248
rect 10296 21188 10300 21244
rect 10300 21188 10356 21244
rect 10356 21188 10360 21244
rect 10296 21184 10360 21188
rect 10376 21244 10440 21248
rect 10376 21188 10380 21244
rect 10380 21188 10436 21244
rect 10436 21188 10440 21244
rect 10376 21184 10440 21188
rect 10456 21244 10520 21248
rect 10456 21188 10460 21244
rect 10460 21188 10516 21244
rect 10516 21188 10520 21244
rect 10456 21184 10520 21188
rect 16216 21244 16280 21248
rect 16216 21188 16220 21244
rect 16220 21188 16276 21244
rect 16276 21188 16280 21244
rect 16216 21184 16280 21188
rect 16296 21244 16360 21248
rect 16296 21188 16300 21244
rect 16300 21188 16356 21244
rect 16356 21188 16360 21244
rect 16296 21184 16360 21188
rect 16376 21244 16440 21248
rect 16376 21188 16380 21244
rect 16380 21188 16436 21244
rect 16436 21188 16440 21244
rect 16376 21184 16440 21188
rect 16456 21244 16520 21248
rect 16456 21188 16460 21244
rect 16460 21188 16516 21244
rect 16516 21188 16520 21244
rect 16456 21184 16520 21188
rect 7216 20700 7280 20704
rect 7216 20644 7220 20700
rect 7220 20644 7276 20700
rect 7276 20644 7280 20700
rect 7216 20640 7280 20644
rect 7296 20700 7360 20704
rect 7296 20644 7300 20700
rect 7300 20644 7356 20700
rect 7356 20644 7360 20700
rect 7296 20640 7360 20644
rect 7376 20700 7440 20704
rect 7376 20644 7380 20700
rect 7380 20644 7436 20700
rect 7436 20644 7440 20700
rect 7376 20640 7440 20644
rect 7456 20700 7520 20704
rect 7456 20644 7460 20700
rect 7460 20644 7516 20700
rect 7516 20644 7520 20700
rect 7456 20640 7520 20644
rect 13216 20700 13280 20704
rect 13216 20644 13220 20700
rect 13220 20644 13276 20700
rect 13276 20644 13280 20700
rect 13216 20640 13280 20644
rect 13296 20700 13360 20704
rect 13296 20644 13300 20700
rect 13300 20644 13356 20700
rect 13356 20644 13360 20700
rect 13296 20640 13360 20644
rect 13376 20700 13440 20704
rect 13376 20644 13380 20700
rect 13380 20644 13436 20700
rect 13436 20644 13440 20700
rect 13376 20640 13440 20644
rect 13456 20700 13520 20704
rect 13456 20644 13460 20700
rect 13460 20644 13516 20700
rect 13516 20644 13520 20700
rect 13456 20640 13520 20644
rect 19216 20700 19280 20704
rect 19216 20644 19220 20700
rect 19220 20644 19276 20700
rect 19276 20644 19280 20700
rect 19216 20640 19280 20644
rect 19296 20700 19360 20704
rect 19296 20644 19300 20700
rect 19300 20644 19356 20700
rect 19356 20644 19360 20700
rect 19296 20640 19360 20644
rect 19376 20700 19440 20704
rect 19376 20644 19380 20700
rect 19380 20644 19436 20700
rect 19436 20644 19440 20700
rect 19376 20640 19440 20644
rect 19456 20700 19520 20704
rect 19456 20644 19460 20700
rect 19460 20644 19516 20700
rect 19516 20644 19520 20700
rect 19456 20640 19520 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 10216 20156 10280 20160
rect 10216 20100 10220 20156
rect 10220 20100 10276 20156
rect 10276 20100 10280 20156
rect 10216 20096 10280 20100
rect 10296 20156 10360 20160
rect 10296 20100 10300 20156
rect 10300 20100 10356 20156
rect 10356 20100 10360 20156
rect 10296 20096 10360 20100
rect 10376 20156 10440 20160
rect 10376 20100 10380 20156
rect 10380 20100 10436 20156
rect 10436 20100 10440 20156
rect 10376 20096 10440 20100
rect 10456 20156 10520 20160
rect 10456 20100 10460 20156
rect 10460 20100 10516 20156
rect 10516 20100 10520 20156
rect 10456 20096 10520 20100
rect 16216 20156 16280 20160
rect 16216 20100 16220 20156
rect 16220 20100 16276 20156
rect 16276 20100 16280 20156
rect 16216 20096 16280 20100
rect 16296 20156 16360 20160
rect 16296 20100 16300 20156
rect 16300 20100 16356 20156
rect 16356 20100 16360 20156
rect 16296 20096 16360 20100
rect 16376 20156 16440 20160
rect 16376 20100 16380 20156
rect 16380 20100 16436 20156
rect 16436 20100 16440 20156
rect 16376 20096 16440 20100
rect 16456 20156 16520 20160
rect 16456 20100 16460 20156
rect 16460 20100 16516 20156
rect 16516 20100 16520 20156
rect 16456 20096 16520 20100
rect 7216 19612 7280 19616
rect 7216 19556 7220 19612
rect 7220 19556 7276 19612
rect 7276 19556 7280 19612
rect 7216 19552 7280 19556
rect 7296 19612 7360 19616
rect 7296 19556 7300 19612
rect 7300 19556 7356 19612
rect 7356 19556 7360 19612
rect 7296 19552 7360 19556
rect 7376 19612 7440 19616
rect 7376 19556 7380 19612
rect 7380 19556 7436 19612
rect 7436 19556 7440 19612
rect 7376 19552 7440 19556
rect 7456 19612 7520 19616
rect 7456 19556 7460 19612
rect 7460 19556 7516 19612
rect 7516 19556 7520 19612
rect 7456 19552 7520 19556
rect 13216 19612 13280 19616
rect 13216 19556 13220 19612
rect 13220 19556 13276 19612
rect 13276 19556 13280 19612
rect 13216 19552 13280 19556
rect 13296 19612 13360 19616
rect 13296 19556 13300 19612
rect 13300 19556 13356 19612
rect 13356 19556 13360 19612
rect 13296 19552 13360 19556
rect 13376 19612 13440 19616
rect 13376 19556 13380 19612
rect 13380 19556 13436 19612
rect 13436 19556 13440 19612
rect 13376 19552 13440 19556
rect 13456 19612 13520 19616
rect 13456 19556 13460 19612
rect 13460 19556 13516 19612
rect 13516 19556 13520 19612
rect 13456 19552 13520 19556
rect 19216 19612 19280 19616
rect 19216 19556 19220 19612
rect 19220 19556 19276 19612
rect 19276 19556 19280 19612
rect 19216 19552 19280 19556
rect 19296 19612 19360 19616
rect 19296 19556 19300 19612
rect 19300 19556 19356 19612
rect 19356 19556 19360 19612
rect 19296 19552 19360 19556
rect 19376 19612 19440 19616
rect 19376 19556 19380 19612
rect 19380 19556 19436 19612
rect 19436 19556 19440 19612
rect 19376 19552 19440 19556
rect 19456 19612 19520 19616
rect 19456 19556 19460 19612
rect 19460 19556 19516 19612
rect 19516 19556 19520 19612
rect 19456 19552 19520 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 10216 19068 10280 19072
rect 10216 19012 10220 19068
rect 10220 19012 10276 19068
rect 10276 19012 10280 19068
rect 10216 19008 10280 19012
rect 10296 19068 10360 19072
rect 10296 19012 10300 19068
rect 10300 19012 10356 19068
rect 10356 19012 10360 19068
rect 10296 19008 10360 19012
rect 10376 19068 10440 19072
rect 10376 19012 10380 19068
rect 10380 19012 10436 19068
rect 10436 19012 10440 19068
rect 10376 19008 10440 19012
rect 10456 19068 10520 19072
rect 10456 19012 10460 19068
rect 10460 19012 10516 19068
rect 10516 19012 10520 19068
rect 10456 19008 10520 19012
rect 16216 19068 16280 19072
rect 16216 19012 16220 19068
rect 16220 19012 16276 19068
rect 16276 19012 16280 19068
rect 16216 19008 16280 19012
rect 16296 19068 16360 19072
rect 16296 19012 16300 19068
rect 16300 19012 16356 19068
rect 16356 19012 16360 19068
rect 16296 19008 16360 19012
rect 16376 19068 16440 19072
rect 16376 19012 16380 19068
rect 16380 19012 16436 19068
rect 16436 19012 16440 19068
rect 16376 19008 16440 19012
rect 16456 19068 16520 19072
rect 16456 19012 16460 19068
rect 16460 19012 16516 19068
rect 16516 19012 16520 19068
rect 16456 19008 16520 19012
rect 7216 18524 7280 18528
rect 7216 18468 7220 18524
rect 7220 18468 7276 18524
rect 7276 18468 7280 18524
rect 7216 18464 7280 18468
rect 7296 18524 7360 18528
rect 7296 18468 7300 18524
rect 7300 18468 7356 18524
rect 7356 18468 7360 18524
rect 7296 18464 7360 18468
rect 7376 18524 7440 18528
rect 7376 18468 7380 18524
rect 7380 18468 7436 18524
rect 7436 18468 7440 18524
rect 7376 18464 7440 18468
rect 7456 18524 7520 18528
rect 7456 18468 7460 18524
rect 7460 18468 7516 18524
rect 7516 18468 7520 18524
rect 7456 18464 7520 18468
rect 13216 18524 13280 18528
rect 13216 18468 13220 18524
rect 13220 18468 13276 18524
rect 13276 18468 13280 18524
rect 13216 18464 13280 18468
rect 13296 18524 13360 18528
rect 13296 18468 13300 18524
rect 13300 18468 13356 18524
rect 13356 18468 13360 18524
rect 13296 18464 13360 18468
rect 13376 18524 13440 18528
rect 13376 18468 13380 18524
rect 13380 18468 13436 18524
rect 13436 18468 13440 18524
rect 13376 18464 13440 18468
rect 13456 18524 13520 18528
rect 13456 18468 13460 18524
rect 13460 18468 13516 18524
rect 13516 18468 13520 18524
rect 13456 18464 13520 18468
rect 19216 18524 19280 18528
rect 19216 18468 19220 18524
rect 19220 18468 19276 18524
rect 19276 18468 19280 18524
rect 19216 18464 19280 18468
rect 19296 18524 19360 18528
rect 19296 18468 19300 18524
rect 19300 18468 19356 18524
rect 19356 18468 19360 18524
rect 19296 18464 19360 18468
rect 19376 18524 19440 18528
rect 19376 18468 19380 18524
rect 19380 18468 19436 18524
rect 19436 18468 19440 18524
rect 19376 18464 19440 18468
rect 19456 18524 19520 18528
rect 19456 18468 19460 18524
rect 19460 18468 19516 18524
rect 19516 18468 19520 18524
rect 19456 18464 19520 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 10216 17980 10280 17984
rect 10216 17924 10220 17980
rect 10220 17924 10276 17980
rect 10276 17924 10280 17980
rect 10216 17920 10280 17924
rect 10296 17980 10360 17984
rect 10296 17924 10300 17980
rect 10300 17924 10356 17980
rect 10356 17924 10360 17980
rect 10296 17920 10360 17924
rect 10376 17980 10440 17984
rect 10376 17924 10380 17980
rect 10380 17924 10436 17980
rect 10436 17924 10440 17980
rect 10376 17920 10440 17924
rect 10456 17980 10520 17984
rect 10456 17924 10460 17980
rect 10460 17924 10516 17980
rect 10516 17924 10520 17980
rect 10456 17920 10520 17924
rect 16216 17980 16280 17984
rect 16216 17924 16220 17980
rect 16220 17924 16276 17980
rect 16276 17924 16280 17980
rect 16216 17920 16280 17924
rect 16296 17980 16360 17984
rect 16296 17924 16300 17980
rect 16300 17924 16356 17980
rect 16356 17924 16360 17980
rect 16296 17920 16360 17924
rect 16376 17980 16440 17984
rect 16376 17924 16380 17980
rect 16380 17924 16436 17980
rect 16436 17924 16440 17980
rect 16376 17920 16440 17924
rect 16456 17980 16520 17984
rect 16456 17924 16460 17980
rect 16460 17924 16516 17980
rect 16516 17924 16520 17980
rect 16456 17920 16520 17924
rect 7216 17436 7280 17440
rect 7216 17380 7220 17436
rect 7220 17380 7276 17436
rect 7276 17380 7280 17436
rect 7216 17376 7280 17380
rect 7296 17436 7360 17440
rect 7296 17380 7300 17436
rect 7300 17380 7356 17436
rect 7356 17380 7360 17436
rect 7296 17376 7360 17380
rect 7376 17436 7440 17440
rect 7376 17380 7380 17436
rect 7380 17380 7436 17436
rect 7436 17380 7440 17436
rect 7376 17376 7440 17380
rect 7456 17436 7520 17440
rect 7456 17380 7460 17436
rect 7460 17380 7516 17436
rect 7516 17380 7520 17436
rect 7456 17376 7520 17380
rect 13216 17436 13280 17440
rect 13216 17380 13220 17436
rect 13220 17380 13276 17436
rect 13276 17380 13280 17436
rect 13216 17376 13280 17380
rect 13296 17436 13360 17440
rect 13296 17380 13300 17436
rect 13300 17380 13356 17436
rect 13356 17380 13360 17436
rect 13296 17376 13360 17380
rect 13376 17436 13440 17440
rect 13376 17380 13380 17436
rect 13380 17380 13436 17436
rect 13436 17380 13440 17436
rect 13376 17376 13440 17380
rect 13456 17436 13520 17440
rect 13456 17380 13460 17436
rect 13460 17380 13516 17436
rect 13516 17380 13520 17436
rect 13456 17376 13520 17380
rect 19216 17436 19280 17440
rect 19216 17380 19220 17436
rect 19220 17380 19276 17436
rect 19276 17380 19280 17436
rect 19216 17376 19280 17380
rect 19296 17436 19360 17440
rect 19296 17380 19300 17436
rect 19300 17380 19356 17436
rect 19356 17380 19360 17436
rect 19296 17376 19360 17380
rect 19376 17436 19440 17440
rect 19376 17380 19380 17436
rect 19380 17380 19436 17436
rect 19436 17380 19440 17436
rect 19376 17376 19440 17380
rect 19456 17436 19520 17440
rect 19456 17380 19460 17436
rect 19460 17380 19516 17436
rect 19516 17380 19520 17436
rect 19456 17376 19520 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 10216 16892 10280 16896
rect 10216 16836 10220 16892
rect 10220 16836 10276 16892
rect 10276 16836 10280 16892
rect 10216 16832 10280 16836
rect 10296 16892 10360 16896
rect 10296 16836 10300 16892
rect 10300 16836 10356 16892
rect 10356 16836 10360 16892
rect 10296 16832 10360 16836
rect 10376 16892 10440 16896
rect 10376 16836 10380 16892
rect 10380 16836 10436 16892
rect 10436 16836 10440 16892
rect 10376 16832 10440 16836
rect 10456 16892 10520 16896
rect 10456 16836 10460 16892
rect 10460 16836 10516 16892
rect 10516 16836 10520 16892
rect 10456 16832 10520 16836
rect 16216 16892 16280 16896
rect 16216 16836 16220 16892
rect 16220 16836 16276 16892
rect 16276 16836 16280 16892
rect 16216 16832 16280 16836
rect 16296 16892 16360 16896
rect 16296 16836 16300 16892
rect 16300 16836 16356 16892
rect 16356 16836 16360 16892
rect 16296 16832 16360 16836
rect 16376 16892 16440 16896
rect 16376 16836 16380 16892
rect 16380 16836 16436 16892
rect 16436 16836 16440 16892
rect 16376 16832 16440 16836
rect 16456 16892 16520 16896
rect 16456 16836 16460 16892
rect 16460 16836 16516 16892
rect 16516 16836 16520 16892
rect 16456 16832 16520 16836
rect 7216 16348 7280 16352
rect 7216 16292 7220 16348
rect 7220 16292 7276 16348
rect 7276 16292 7280 16348
rect 7216 16288 7280 16292
rect 7296 16348 7360 16352
rect 7296 16292 7300 16348
rect 7300 16292 7356 16348
rect 7356 16292 7360 16348
rect 7296 16288 7360 16292
rect 7376 16348 7440 16352
rect 7376 16292 7380 16348
rect 7380 16292 7436 16348
rect 7436 16292 7440 16348
rect 7376 16288 7440 16292
rect 7456 16348 7520 16352
rect 7456 16292 7460 16348
rect 7460 16292 7516 16348
rect 7516 16292 7520 16348
rect 7456 16288 7520 16292
rect 13216 16348 13280 16352
rect 13216 16292 13220 16348
rect 13220 16292 13276 16348
rect 13276 16292 13280 16348
rect 13216 16288 13280 16292
rect 13296 16348 13360 16352
rect 13296 16292 13300 16348
rect 13300 16292 13356 16348
rect 13356 16292 13360 16348
rect 13296 16288 13360 16292
rect 13376 16348 13440 16352
rect 13376 16292 13380 16348
rect 13380 16292 13436 16348
rect 13436 16292 13440 16348
rect 13376 16288 13440 16292
rect 13456 16348 13520 16352
rect 13456 16292 13460 16348
rect 13460 16292 13516 16348
rect 13516 16292 13520 16348
rect 13456 16288 13520 16292
rect 19216 16348 19280 16352
rect 19216 16292 19220 16348
rect 19220 16292 19276 16348
rect 19276 16292 19280 16348
rect 19216 16288 19280 16292
rect 19296 16348 19360 16352
rect 19296 16292 19300 16348
rect 19300 16292 19356 16348
rect 19356 16292 19360 16348
rect 19296 16288 19360 16292
rect 19376 16348 19440 16352
rect 19376 16292 19380 16348
rect 19380 16292 19436 16348
rect 19436 16292 19440 16348
rect 19376 16288 19440 16292
rect 19456 16348 19520 16352
rect 19456 16292 19460 16348
rect 19460 16292 19516 16348
rect 19516 16292 19520 16348
rect 19456 16288 19520 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 10216 15804 10280 15808
rect 10216 15748 10220 15804
rect 10220 15748 10276 15804
rect 10276 15748 10280 15804
rect 10216 15744 10280 15748
rect 10296 15804 10360 15808
rect 10296 15748 10300 15804
rect 10300 15748 10356 15804
rect 10356 15748 10360 15804
rect 10296 15744 10360 15748
rect 10376 15804 10440 15808
rect 10376 15748 10380 15804
rect 10380 15748 10436 15804
rect 10436 15748 10440 15804
rect 10376 15744 10440 15748
rect 10456 15804 10520 15808
rect 10456 15748 10460 15804
rect 10460 15748 10516 15804
rect 10516 15748 10520 15804
rect 10456 15744 10520 15748
rect 16216 15804 16280 15808
rect 16216 15748 16220 15804
rect 16220 15748 16276 15804
rect 16276 15748 16280 15804
rect 16216 15744 16280 15748
rect 16296 15804 16360 15808
rect 16296 15748 16300 15804
rect 16300 15748 16356 15804
rect 16356 15748 16360 15804
rect 16296 15744 16360 15748
rect 16376 15804 16440 15808
rect 16376 15748 16380 15804
rect 16380 15748 16436 15804
rect 16436 15748 16440 15804
rect 16376 15744 16440 15748
rect 16456 15804 16520 15808
rect 16456 15748 16460 15804
rect 16460 15748 16516 15804
rect 16516 15748 16520 15804
rect 16456 15744 16520 15748
rect 7216 15260 7280 15264
rect 7216 15204 7220 15260
rect 7220 15204 7276 15260
rect 7276 15204 7280 15260
rect 7216 15200 7280 15204
rect 7296 15260 7360 15264
rect 7296 15204 7300 15260
rect 7300 15204 7356 15260
rect 7356 15204 7360 15260
rect 7296 15200 7360 15204
rect 7376 15260 7440 15264
rect 7376 15204 7380 15260
rect 7380 15204 7436 15260
rect 7436 15204 7440 15260
rect 7376 15200 7440 15204
rect 7456 15260 7520 15264
rect 7456 15204 7460 15260
rect 7460 15204 7516 15260
rect 7516 15204 7520 15260
rect 7456 15200 7520 15204
rect 13216 15260 13280 15264
rect 13216 15204 13220 15260
rect 13220 15204 13276 15260
rect 13276 15204 13280 15260
rect 13216 15200 13280 15204
rect 13296 15260 13360 15264
rect 13296 15204 13300 15260
rect 13300 15204 13356 15260
rect 13356 15204 13360 15260
rect 13296 15200 13360 15204
rect 13376 15260 13440 15264
rect 13376 15204 13380 15260
rect 13380 15204 13436 15260
rect 13436 15204 13440 15260
rect 13376 15200 13440 15204
rect 13456 15260 13520 15264
rect 13456 15204 13460 15260
rect 13460 15204 13516 15260
rect 13516 15204 13520 15260
rect 13456 15200 13520 15204
rect 19216 15260 19280 15264
rect 19216 15204 19220 15260
rect 19220 15204 19276 15260
rect 19276 15204 19280 15260
rect 19216 15200 19280 15204
rect 19296 15260 19360 15264
rect 19296 15204 19300 15260
rect 19300 15204 19356 15260
rect 19356 15204 19360 15260
rect 19296 15200 19360 15204
rect 19376 15260 19440 15264
rect 19376 15204 19380 15260
rect 19380 15204 19436 15260
rect 19436 15204 19440 15260
rect 19376 15200 19440 15204
rect 19456 15260 19520 15264
rect 19456 15204 19460 15260
rect 19460 15204 19516 15260
rect 19516 15204 19520 15260
rect 19456 15200 19520 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 10216 14716 10280 14720
rect 10216 14660 10220 14716
rect 10220 14660 10276 14716
rect 10276 14660 10280 14716
rect 10216 14656 10280 14660
rect 10296 14716 10360 14720
rect 10296 14660 10300 14716
rect 10300 14660 10356 14716
rect 10356 14660 10360 14716
rect 10296 14656 10360 14660
rect 10376 14716 10440 14720
rect 10376 14660 10380 14716
rect 10380 14660 10436 14716
rect 10436 14660 10440 14716
rect 10376 14656 10440 14660
rect 10456 14716 10520 14720
rect 10456 14660 10460 14716
rect 10460 14660 10516 14716
rect 10516 14660 10520 14716
rect 10456 14656 10520 14660
rect 16216 14716 16280 14720
rect 16216 14660 16220 14716
rect 16220 14660 16276 14716
rect 16276 14660 16280 14716
rect 16216 14656 16280 14660
rect 16296 14716 16360 14720
rect 16296 14660 16300 14716
rect 16300 14660 16356 14716
rect 16356 14660 16360 14716
rect 16296 14656 16360 14660
rect 16376 14716 16440 14720
rect 16376 14660 16380 14716
rect 16380 14660 16436 14716
rect 16436 14660 16440 14716
rect 16376 14656 16440 14660
rect 16456 14716 16520 14720
rect 16456 14660 16460 14716
rect 16460 14660 16516 14716
rect 16516 14660 16520 14716
rect 16456 14656 16520 14660
rect 7216 14172 7280 14176
rect 7216 14116 7220 14172
rect 7220 14116 7276 14172
rect 7276 14116 7280 14172
rect 7216 14112 7280 14116
rect 7296 14172 7360 14176
rect 7296 14116 7300 14172
rect 7300 14116 7356 14172
rect 7356 14116 7360 14172
rect 7296 14112 7360 14116
rect 7376 14172 7440 14176
rect 7376 14116 7380 14172
rect 7380 14116 7436 14172
rect 7436 14116 7440 14172
rect 7376 14112 7440 14116
rect 7456 14172 7520 14176
rect 7456 14116 7460 14172
rect 7460 14116 7516 14172
rect 7516 14116 7520 14172
rect 7456 14112 7520 14116
rect 13216 14172 13280 14176
rect 13216 14116 13220 14172
rect 13220 14116 13276 14172
rect 13276 14116 13280 14172
rect 13216 14112 13280 14116
rect 13296 14172 13360 14176
rect 13296 14116 13300 14172
rect 13300 14116 13356 14172
rect 13356 14116 13360 14172
rect 13296 14112 13360 14116
rect 13376 14172 13440 14176
rect 13376 14116 13380 14172
rect 13380 14116 13436 14172
rect 13436 14116 13440 14172
rect 13376 14112 13440 14116
rect 13456 14172 13520 14176
rect 13456 14116 13460 14172
rect 13460 14116 13516 14172
rect 13516 14116 13520 14172
rect 13456 14112 13520 14116
rect 19216 14172 19280 14176
rect 19216 14116 19220 14172
rect 19220 14116 19276 14172
rect 19276 14116 19280 14172
rect 19216 14112 19280 14116
rect 19296 14172 19360 14176
rect 19296 14116 19300 14172
rect 19300 14116 19356 14172
rect 19356 14116 19360 14172
rect 19296 14112 19360 14116
rect 19376 14172 19440 14176
rect 19376 14116 19380 14172
rect 19380 14116 19436 14172
rect 19436 14116 19440 14172
rect 19376 14112 19440 14116
rect 19456 14172 19520 14176
rect 19456 14116 19460 14172
rect 19460 14116 19516 14172
rect 19516 14116 19520 14172
rect 19456 14112 19520 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 10216 13628 10280 13632
rect 10216 13572 10220 13628
rect 10220 13572 10276 13628
rect 10276 13572 10280 13628
rect 10216 13568 10280 13572
rect 10296 13628 10360 13632
rect 10296 13572 10300 13628
rect 10300 13572 10356 13628
rect 10356 13572 10360 13628
rect 10296 13568 10360 13572
rect 10376 13628 10440 13632
rect 10376 13572 10380 13628
rect 10380 13572 10436 13628
rect 10436 13572 10440 13628
rect 10376 13568 10440 13572
rect 10456 13628 10520 13632
rect 10456 13572 10460 13628
rect 10460 13572 10516 13628
rect 10516 13572 10520 13628
rect 10456 13568 10520 13572
rect 16216 13628 16280 13632
rect 16216 13572 16220 13628
rect 16220 13572 16276 13628
rect 16276 13572 16280 13628
rect 16216 13568 16280 13572
rect 16296 13628 16360 13632
rect 16296 13572 16300 13628
rect 16300 13572 16356 13628
rect 16356 13572 16360 13628
rect 16296 13568 16360 13572
rect 16376 13628 16440 13632
rect 16376 13572 16380 13628
rect 16380 13572 16436 13628
rect 16436 13572 16440 13628
rect 16376 13568 16440 13572
rect 16456 13628 16520 13632
rect 16456 13572 16460 13628
rect 16460 13572 16516 13628
rect 16516 13572 16520 13628
rect 16456 13568 16520 13572
rect 7216 13084 7280 13088
rect 7216 13028 7220 13084
rect 7220 13028 7276 13084
rect 7276 13028 7280 13084
rect 7216 13024 7280 13028
rect 7296 13084 7360 13088
rect 7296 13028 7300 13084
rect 7300 13028 7356 13084
rect 7356 13028 7360 13084
rect 7296 13024 7360 13028
rect 7376 13084 7440 13088
rect 7376 13028 7380 13084
rect 7380 13028 7436 13084
rect 7436 13028 7440 13084
rect 7376 13024 7440 13028
rect 7456 13084 7520 13088
rect 7456 13028 7460 13084
rect 7460 13028 7516 13084
rect 7516 13028 7520 13084
rect 7456 13024 7520 13028
rect 13216 13084 13280 13088
rect 13216 13028 13220 13084
rect 13220 13028 13276 13084
rect 13276 13028 13280 13084
rect 13216 13024 13280 13028
rect 13296 13084 13360 13088
rect 13296 13028 13300 13084
rect 13300 13028 13356 13084
rect 13356 13028 13360 13084
rect 13296 13024 13360 13028
rect 13376 13084 13440 13088
rect 13376 13028 13380 13084
rect 13380 13028 13436 13084
rect 13436 13028 13440 13084
rect 13376 13024 13440 13028
rect 13456 13084 13520 13088
rect 13456 13028 13460 13084
rect 13460 13028 13516 13084
rect 13516 13028 13520 13084
rect 13456 13024 13520 13028
rect 19216 13084 19280 13088
rect 19216 13028 19220 13084
rect 19220 13028 19276 13084
rect 19276 13028 19280 13084
rect 19216 13024 19280 13028
rect 19296 13084 19360 13088
rect 19296 13028 19300 13084
rect 19300 13028 19356 13084
rect 19356 13028 19360 13084
rect 19296 13024 19360 13028
rect 19376 13084 19440 13088
rect 19376 13028 19380 13084
rect 19380 13028 19436 13084
rect 19436 13028 19440 13084
rect 19376 13024 19440 13028
rect 19456 13084 19520 13088
rect 19456 13028 19460 13084
rect 19460 13028 19516 13084
rect 19516 13028 19520 13084
rect 19456 13024 19520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 10216 12540 10280 12544
rect 10216 12484 10220 12540
rect 10220 12484 10276 12540
rect 10276 12484 10280 12540
rect 10216 12480 10280 12484
rect 10296 12540 10360 12544
rect 10296 12484 10300 12540
rect 10300 12484 10356 12540
rect 10356 12484 10360 12540
rect 10296 12480 10360 12484
rect 10376 12540 10440 12544
rect 10376 12484 10380 12540
rect 10380 12484 10436 12540
rect 10436 12484 10440 12540
rect 10376 12480 10440 12484
rect 10456 12540 10520 12544
rect 10456 12484 10460 12540
rect 10460 12484 10516 12540
rect 10516 12484 10520 12540
rect 10456 12480 10520 12484
rect 16216 12540 16280 12544
rect 16216 12484 16220 12540
rect 16220 12484 16276 12540
rect 16276 12484 16280 12540
rect 16216 12480 16280 12484
rect 16296 12540 16360 12544
rect 16296 12484 16300 12540
rect 16300 12484 16356 12540
rect 16356 12484 16360 12540
rect 16296 12480 16360 12484
rect 16376 12540 16440 12544
rect 16376 12484 16380 12540
rect 16380 12484 16436 12540
rect 16436 12484 16440 12540
rect 16376 12480 16440 12484
rect 16456 12540 16520 12544
rect 16456 12484 16460 12540
rect 16460 12484 16516 12540
rect 16516 12484 16520 12540
rect 16456 12480 16520 12484
rect 7216 11996 7280 12000
rect 7216 11940 7220 11996
rect 7220 11940 7276 11996
rect 7276 11940 7280 11996
rect 7216 11936 7280 11940
rect 7296 11996 7360 12000
rect 7296 11940 7300 11996
rect 7300 11940 7356 11996
rect 7356 11940 7360 11996
rect 7296 11936 7360 11940
rect 7376 11996 7440 12000
rect 7376 11940 7380 11996
rect 7380 11940 7436 11996
rect 7436 11940 7440 11996
rect 7376 11936 7440 11940
rect 7456 11996 7520 12000
rect 7456 11940 7460 11996
rect 7460 11940 7516 11996
rect 7516 11940 7520 11996
rect 7456 11936 7520 11940
rect 13216 11996 13280 12000
rect 13216 11940 13220 11996
rect 13220 11940 13276 11996
rect 13276 11940 13280 11996
rect 13216 11936 13280 11940
rect 13296 11996 13360 12000
rect 13296 11940 13300 11996
rect 13300 11940 13356 11996
rect 13356 11940 13360 11996
rect 13296 11936 13360 11940
rect 13376 11996 13440 12000
rect 13376 11940 13380 11996
rect 13380 11940 13436 11996
rect 13436 11940 13440 11996
rect 13376 11936 13440 11940
rect 13456 11996 13520 12000
rect 13456 11940 13460 11996
rect 13460 11940 13516 11996
rect 13516 11940 13520 11996
rect 13456 11936 13520 11940
rect 19216 11996 19280 12000
rect 19216 11940 19220 11996
rect 19220 11940 19276 11996
rect 19276 11940 19280 11996
rect 19216 11936 19280 11940
rect 19296 11996 19360 12000
rect 19296 11940 19300 11996
rect 19300 11940 19356 11996
rect 19356 11940 19360 11996
rect 19296 11936 19360 11940
rect 19376 11996 19440 12000
rect 19376 11940 19380 11996
rect 19380 11940 19436 11996
rect 19436 11940 19440 11996
rect 19376 11936 19440 11940
rect 19456 11996 19520 12000
rect 19456 11940 19460 11996
rect 19460 11940 19516 11996
rect 19516 11940 19520 11996
rect 19456 11936 19520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 10216 11452 10280 11456
rect 10216 11396 10220 11452
rect 10220 11396 10276 11452
rect 10276 11396 10280 11452
rect 10216 11392 10280 11396
rect 10296 11452 10360 11456
rect 10296 11396 10300 11452
rect 10300 11396 10356 11452
rect 10356 11396 10360 11452
rect 10296 11392 10360 11396
rect 10376 11452 10440 11456
rect 10376 11396 10380 11452
rect 10380 11396 10436 11452
rect 10436 11396 10440 11452
rect 10376 11392 10440 11396
rect 10456 11452 10520 11456
rect 10456 11396 10460 11452
rect 10460 11396 10516 11452
rect 10516 11396 10520 11452
rect 10456 11392 10520 11396
rect 16216 11452 16280 11456
rect 16216 11396 16220 11452
rect 16220 11396 16276 11452
rect 16276 11396 16280 11452
rect 16216 11392 16280 11396
rect 16296 11452 16360 11456
rect 16296 11396 16300 11452
rect 16300 11396 16356 11452
rect 16356 11396 16360 11452
rect 16296 11392 16360 11396
rect 16376 11452 16440 11456
rect 16376 11396 16380 11452
rect 16380 11396 16436 11452
rect 16436 11396 16440 11452
rect 16376 11392 16440 11396
rect 16456 11452 16520 11456
rect 16456 11396 16460 11452
rect 16460 11396 16516 11452
rect 16516 11396 16520 11452
rect 16456 11392 16520 11396
rect 7216 10908 7280 10912
rect 7216 10852 7220 10908
rect 7220 10852 7276 10908
rect 7276 10852 7280 10908
rect 7216 10848 7280 10852
rect 7296 10908 7360 10912
rect 7296 10852 7300 10908
rect 7300 10852 7356 10908
rect 7356 10852 7360 10908
rect 7296 10848 7360 10852
rect 7376 10908 7440 10912
rect 7376 10852 7380 10908
rect 7380 10852 7436 10908
rect 7436 10852 7440 10908
rect 7376 10848 7440 10852
rect 7456 10908 7520 10912
rect 7456 10852 7460 10908
rect 7460 10852 7516 10908
rect 7516 10852 7520 10908
rect 7456 10848 7520 10852
rect 13216 10908 13280 10912
rect 13216 10852 13220 10908
rect 13220 10852 13276 10908
rect 13276 10852 13280 10908
rect 13216 10848 13280 10852
rect 13296 10908 13360 10912
rect 13296 10852 13300 10908
rect 13300 10852 13356 10908
rect 13356 10852 13360 10908
rect 13296 10848 13360 10852
rect 13376 10908 13440 10912
rect 13376 10852 13380 10908
rect 13380 10852 13436 10908
rect 13436 10852 13440 10908
rect 13376 10848 13440 10852
rect 13456 10908 13520 10912
rect 13456 10852 13460 10908
rect 13460 10852 13516 10908
rect 13516 10852 13520 10908
rect 13456 10848 13520 10852
rect 19216 10908 19280 10912
rect 19216 10852 19220 10908
rect 19220 10852 19276 10908
rect 19276 10852 19280 10908
rect 19216 10848 19280 10852
rect 19296 10908 19360 10912
rect 19296 10852 19300 10908
rect 19300 10852 19356 10908
rect 19356 10852 19360 10908
rect 19296 10848 19360 10852
rect 19376 10908 19440 10912
rect 19376 10852 19380 10908
rect 19380 10852 19436 10908
rect 19436 10852 19440 10908
rect 19376 10848 19440 10852
rect 19456 10908 19520 10912
rect 19456 10852 19460 10908
rect 19460 10852 19516 10908
rect 19516 10852 19520 10908
rect 19456 10848 19520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 10216 10364 10280 10368
rect 10216 10308 10220 10364
rect 10220 10308 10276 10364
rect 10276 10308 10280 10364
rect 10216 10304 10280 10308
rect 10296 10364 10360 10368
rect 10296 10308 10300 10364
rect 10300 10308 10356 10364
rect 10356 10308 10360 10364
rect 10296 10304 10360 10308
rect 10376 10364 10440 10368
rect 10376 10308 10380 10364
rect 10380 10308 10436 10364
rect 10436 10308 10440 10364
rect 10376 10304 10440 10308
rect 10456 10364 10520 10368
rect 10456 10308 10460 10364
rect 10460 10308 10516 10364
rect 10516 10308 10520 10364
rect 10456 10304 10520 10308
rect 16216 10364 16280 10368
rect 16216 10308 16220 10364
rect 16220 10308 16276 10364
rect 16276 10308 16280 10364
rect 16216 10304 16280 10308
rect 16296 10364 16360 10368
rect 16296 10308 16300 10364
rect 16300 10308 16356 10364
rect 16356 10308 16360 10364
rect 16296 10304 16360 10308
rect 16376 10364 16440 10368
rect 16376 10308 16380 10364
rect 16380 10308 16436 10364
rect 16436 10308 16440 10364
rect 16376 10304 16440 10308
rect 16456 10364 16520 10368
rect 16456 10308 16460 10364
rect 16460 10308 16516 10364
rect 16516 10308 16520 10364
rect 16456 10304 16520 10308
rect 7216 9820 7280 9824
rect 7216 9764 7220 9820
rect 7220 9764 7276 9820
rect 7276 9764 7280 9820
rect 7216 9760 7280 9764
rect 7296 9820 7360 9824
rect 7296 9764 7300 9820
rect 7300 9764 7356 9820
rect 7356 9764 7360 9820
rect 7296 9760 7360 9764
rect 7376 9820 7440 9824
rect 7376 9764 7380 9820
rect 7380 9764 7436 9820
rect 7436 9764 7440 9820
rect 7376 9760 7440 9764
rect 7456 9820 7520 9824
rect 7456 9764 7460 9820
rect 7460 9764 7516 9820
rect 7516 9764 7520 9820
rect 7456 9760 7520 9764
rect 13216 9820 13280 9824
rect 13216 9764 13220 9820
rect 13220 9764 13276 9820
rect 13276 9764 13280 9820
rect 13216 9760 13280 9764
rect 13296 9820 13360 9824
rect 13296 9764 13300 9820
rect 13300 9764 13356 9820
rect 13356 9764 13360 9820
rect 13296 9760 13360 9764
rect 13376 9820 13440 9824
rect 13376 9764 13380 9820
rect 13380 9764 13436 9820
rect 13436 9764 13440 9820
rect 13376 9760 13440 9764
rect 13456 9820 13520 9824
rect 13456 9764 13460 9820
rect 13460 9764 13516 9820
rect 13516 9764 13520 9820
rect 13456 9760 13520 9764
rect 19216 9820 19280 9824
rect 19216 9764 19220 9820
rect 19220 9764 19276 9820
rect 19276 9764 19280 9820
rect 19216 9760 19280 9764
rect 19296 9820 19360 9824
rect 19296 9764 19300 9820
rect 19300 9764 19356 9820
rect 19356 9764 19360 9820
rect 19296 9760 19360 9764
rect 19376 9820 19440 9824
rect 19376 9764 19380 9820
rect 19380 9764 19436 9820
rect 19436 9764 19440 9820
rect 19376 9760 19440 9764
rect 19456 9820 19520 9824
rect 19456 9764 19460 9820
rect 19460 9764 19516 9820
rect 19516 9764 19520 9820
rect 19456 9760 19520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 10216 9276 10280 9280
rect 10216 9220 10220 9276
rect 10220 9220 10276 9276
rect 10276 9220 10280 9276
rect 10216 9216 10280 9220
rect 10296 9276 10360 9280
rect 10296 9220 10300 9276
rect 10300 9220 10356 9276
rect 10356 9220 10360 9276
rect 10296 9216 10360 9220
rect 10376 9276 10440 9280
rect 10376 9220 10380 9276
rect 10380 9220 10436 9276
rect 10436 9220 10440 9276
rect 10376 9216 10440 9220
rect 10456 9276 10520 9280
rect 10456 9220 10460 9276
rect 10460 9220 10516 9276
rect 10516 9220 10520 9276
rect 10456 9216 10520 9220
rect 16216 9276 16280 9280
rect 16216 9220 16220 9276
rect 16220 9220 16276 9276
rect 16276 9220 16280 9276
rect 16216 9216 16280 9220
rect 16296 9276 16360 9280
rect 16296 9220 16300 9276
rect 16300 9220 16356 9276
rect 16356 9220 16360 9276
rect 16296 9216 16360 9220
rect 16376 9276 16440 9280
rect 16376 9220 16380 9276
rect 16380 9220 16436 9276
rect 16436 9220 16440 9276
rect 16376 9216 16440 9220
rect 16456 9276 16520 9280
rect 16456 9220 16460 9276
rect 16460 9220 16516 9276
rect 16516 9220 16520 9276
rect 16456 9216 16520 9220
rect 7216 8732 7280 8736
rect 7216 8676 7220 8732
rect 7220 8676 7276 8732
rect 7276 8676 7280 8732
rect 7216 8672 7280 8676
rect 7296 8732 7360 8736
rect 7296 8676 7300 8732
rect 7300 8676 7356 8732
rect 7356 8676 7360 8732
rect 7296 8672 7360 8676
rect 7376 8732 7440 8736
rect 7376 8676 7380 8732
rect 7380 8676 7436 8732
rect 7436 8676 7440 8732
rect 7376 8672 7440 8676
rect 7456 8732 7520 8736
rect 7456 8676 7460 8732
rect 7460 8676 7516 8732
rect 7516 8676 7520 8732
rect 7456 8672 7520 8676
rect 13216 8732 13280 8736
rect 13216 8676 13220 8732
rect 13220 8676 13276 8732
rect 13276 8676 13280 8732
rect 13216 8672 13280 8676
rect 13296 8732 13360 8736
rect 13296 8676 13300 8732
rect 13300 8676 13356 8732
rect 13356 8676 13360 8732
rect 13296 8672 13360 8676
rect 13376 8732 13440 8736
rect 13376 8676 13380 8732
rect 13380 8676 13436 8732
rect 13436 8676 13440 8732
rect 13376 8672 13440 8676
rect 13456 8732 13520 8736
rect 13456 8676 13460 8732
rect 13460 8676 13516 8732
rect 13516 8676 13520 8732
rect 13456 8672 13520 8676
rect 19216 8732 19280 8736
rect 19216 8676 19220 8732
rect 19220 8676 19276 8732
rect 19276 8676 19280 8732
rect 19216 8672 19280 8676
rect 19296 8732 19360 8736
rect 19296 8676 19300 8732
rect 19300 8676 19356 8732
rect 19356 8676 19360 8732
rect 19296 8672 19360 8676
rect 19376 8732 19440 8736
rect 19376 8676 19380 8732
rect 19380 8676 19436 8732
rect 19436 8676 19440 8732
rect 19376 8672 19440 8676
rect 19456 8732 19520 8736
rect 19456 8676 19460 8732
rect 19460 8676 19516 8732
rect 19516 8676 19520 8732
rect 19456 8672 19520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 10216 8188 10280 8192
rect 10216 8132 10220 8188
rect 10220 8132 10276 8188
rect 10276 8132 10280 8188
rect 10216 8128 10280 8132
rect 10296 8188 10360 8192
rect 10296 8132 10300 8188
rect 10300 8132 10356 8188
rect 10356 8132 10360 8188
rect 10296 8128 10360 8132
rect 10376 8188 10440 8192
rect 10376 8132 10380 8188
rect 10380 8132 10436 8188
rect 10436 8132 10440 8188
rect 10376 8128 10440 8132
rect 10456 8188 10520 8192
rect 10456 8132 10460 8188
rect 10460 8132 10516 8188
rect 10516 8132 10520 8188
rect 10456 8128 10520 8132
rect 16216 8188 16280 8192
rect 16216 8132 16220 8188
rect 16220 8132 16276 8188
rect 16276 8132 16280 8188
rect 16216 8128 16280 8132
rect 16296 8188 16360 8192
rect 16296 8132 16300 8188
rect 16300 8132 16356 8188
rect 16356 8132 16360 8188
rect 16296 8128 16360 8132
rect 16376 8188 16440 8192
rect 16376 8132 16380 8188
rect 16380 8132 16436 8188
rect 16436 8132 16440 8188
rect 16376 8128 16440 8132
rect 16456 8188 16520 8192
rect 16456 8132 16460 8188
rect 16460 8132 16516 8188
rect 16516 8132 16520 8188
rect 16456 8128 16520 8132
rect 7216 7644 7280 7648
rect 7216 7588 7220 7644
rect 7220 7588 7276 7644
rect 7276 7588 7280 7644
rect 7216 7584 7280 7588
rect 7296 7644 7360 7648
rect 7296 7588 7300 7644
rect 7300 7588 7356 7644
rect 7356 7588 7360 7644
rect 7296 7584 7360 7588
rect 7376 7644 7440 7648
rect 7376 7588 7380 7644
rect 7380 7588 7436 7644
rect 7436 7588 7440 7644
rect 7376 7584 7440 7588
rect 7456 7644 7520 7648
rect 7456 7588 7460 7644
rect 7460 7588 7516 7644
rect 7516 7588 7520 7644
rect 7456 7584 7520 7588
rect 13216 7644 13280 7648
rect 13216 7588 13220 7644
rect 13220 7588 13276 7644
rect 13276 7588 13280 7644
rect 13216 7584 13280 7588
rect 13296 7644 13360 7648
rect 13296 7588 13300 7644
rect 13300 7588 13356 7644
rect 13356 7588 13360 7644
rect 13296 7584 13360 7588
rect 13376 7644 13440 7648
rect 13376 7588 13380 7644
rect 13380 7588 13436 7644
rect 13436 7588 13440 7644
rect 13376 7584 13440 7588
rect 13456 7644 13520 7648
rect 13456 7588 13460 7644
rect 13460 7588 13516 7644
rect 13516 7588 13520 7644
rect 13456 7584 13520 7588
rect 19216 7644 19280 7648
rect 19216 7588 19220 7644
rect 19220 7588 19276 7644
rect 19276 7588 19280 7644
rect 19216 7584 19280 7588
rect 19296 7644 19360 7648
rect 19296 7588 19300 7644
rect 19300 7588 19356 7644
rect 19356 7588 19360 7644
rect 19296 7584 19360 7588
rect 19376 7644 19440 7648
rect 19376 7588 19380 7644
rect 19380 7588 19436 7644
rect 19436 7588 19440 7644
rect 19376 7584 19440 7588
rect 19456 7644 19520 7648
rect 19456 7588 19460 7644
rect 19460 7588 19516 7644
rect 19516 7588 19520 7644
rect 19456 7584 19520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 10216 7100 10280 7104
rect 10216 7044 10220 7100
rect 10220 7044 10276 7100
rect 10276 7044 10280 7100
rect 10216 7040 10280 7044
rect 10296 7100 10360 7104
rect 10296 7044 10300 7100
rect 10300 7044 10356 7100
rect 10356 7044 10360 7100
rect 10296 7040 10360 7044
rect 10376 7100 10440 7104
rect 10376 7044 10380 7100
rect 10380 7044 10436 7100
rect 10436 7044 10440 7100
rect 10376 7040 10440 7044
rect 10456 7100 10520 7104
rect 10456 7044 10460 7100
rect 10460 7044 10516 7100
rect 10516 7044 10520 7100
rect 10456 7040 10520 7044
rect 16216 7100 16280 7104
rect 16216 7044 16220 7100
rect 16220 7044 16276 7100
rect 16276 7044 16280 7100
rect 16216 7040 16280 7044
rect 16296 7100 16360 7104
rect 16296 7044 16300 7100
rect 16300 7044 16356 7100
rect 16356 7044 16360 7100
rect 16296 7040 16360 7044
rect 16376 7100 16440 7104
rect 16376 7044 16380 7100
rect 16380 7044 16436 7100
rect 16436 7044 16440 7100
rect 16376 7040 16440 7044
rect 16456 7100 16520 7104
rect 16456 7044 16460 7100
rect 16460 7044 16516 7100
rect 16516 7044 16520 7100
rect 16456 7040 16520 7044
rect 7216 6556 7280 6560
rect 7216 6500 7220 6556
rect 7220 6500 7276 6556
rect 7276 6500 7280 6556
rect 7216 6496 7280 6500
rect 7296 6556 7360 6560
rect 7296 6500 7300 6556
rect 7300 6500 7356 6556
rect 7356 6500 7360 6556
rect 7296 6496 7360 6500
rect 7376 6556 7440 6560
rect 7376 6500 7380 6556
rect 7380 6500 7436 6556
rect 7436 6500 7440 6556
rect 7376 6496 7440 6500
rect 7456 6556 7520 6560
rect 7456 6500 7460 6556
rect 7460 6500 7516 6556
rect 7516 6500 7520 6556
rect 7456 6496 7520 6500
rect 13216 6556 13280 6560
rect 13216 6500 13220 6556
rect 13220 6500 13276 6556
rect 13276 6500 13280 6556
rect 13216 6496 13280 6500
rect 13296 6556 13360 6560
rect 13296 6500 13300 6556
rect 13300 6500 13356 6556
rect 13356 6500 13360 6556
rect 13296 6496 13360 6500
rect 13376 6556 13440 6560
rect 13376 6500 13380 6556
rect 13380 6500 13436 6556
rect 13436 6500 13440 6556
rect 13376 6496 13440 6500
rect 13456 6556 13520 6560
rect 13456 6500 13460 6556
rect 13460 6500 13516 6556
rect 13516 6500 13520 6556
rect 13456 6496 13520 6500
rect 19216 6556 19280 6560
rect 19216 6500 19220 6556
rect 19220 6500 19276 6556
rect 19276 6500 19280 6556
rect 19216 6496 19280 6500
rect 19296 6556 19360 6560
rect 19296 6500 19300 6556
rect 19300 6500 19356 6556
rect 19356 6500 19360 6556
rect 19296 6496 19360 6500
rect 19376 6556 19440 6560
rect 19376 6500 19380 6556
rect 19380 6500 19436 6556
rect 19436 6500 19440 6556
rect 19376 6496 19440 6500
rect 19456 6556 19520 6560
rect 19456 6500 19460 6556
rect 19460 6500 19516 6556
rect 19516 6500 19520 6556
rect 19456 6496 19520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 10216 6012 10280 6016
rect 10216 5956 10220 6012
rect 10220 5956 10276 6012
rect 10276 5956 10280 6012
rect 10216 5952 10280 5956
rect 10296 6012 10360 6016
rect 10296 5956 10300 6012
rect 10300 5956 10356 6012
rect 10356 5956 10360 6012
rect 10296 5952 10360 5956
rect 10376 6012 10440 6016
rect 10376 5956 10380 6012
rect 10380 5956 10436 6012
rect 10436 5956 10440 6012
rect 10376 5952 10440 5956
rect 10456 6012 10520 6016
rect 10456 5956 10460 6012
rect 10460 5956 10516 6012
rect 10516 5956 10520 6012
rect 10456 5952 10520 5956
rect 16216 6012 16280 6016
rect 16216 5956 16220 6012
rect 16220 5956 16276 6012
rect 16276 5956 16280 6012
rect 16216 5952 16280 5956
rect 16296 6012 16360 6016
rect 16296 5956 16300 6012
rect 16300 5956 16356 6012
rect 16356 5956 16360 6012
rect 16296 5952 16360 5956
rect 16376 6012 16440 6016
rect 16376 5956 16380 6012
rect 16380 5956 16436 6012
rect 16436 5956 16440 6012
rect 16376 5952 16440 5956
rect 16456 6012 16520 6016
rect 16456 5956 16460 6012
rect 16460 5956 16516 6012
rect 16516 5956 16520 6012
rect 16456 5952 16520 5956
rect 7216 5468 7280 5472
rect 7216 5412 7220 5468
rect 7220 5412 7276 5468
rect 7276 5412 7280 5468
rect 7216 5408 7280 5412
rect 7296 5468 7360 5472
rect 7296 5412 7300 5468
rect 7300 5412 7356 5468
rect 7356 5412 7360 5468
rect 7296 5408 7360 5412
rect 7376 5468 7440 5472
rect 7376 5412 7380 5468
rect 7380 5412 7436 5468
rect 7436 5412 7440 5468
rect 7376 5408 7440 5412
rect 7456 5468 7520 5472
rect 7456 5412 7460 5468
rect 7460 5412 7516 5468
rect 7516 5412 7520 5468
rect 7456 5408 7520 5412
rect 13216 5468 13280 5472
rect 13216 5412 13220 5468
rect 13220 5412 13276 5468
rect 13276 5412 13280 5468
rect 13216 5408 13280 5412
rect 13296 5468 13360 5472
rect 13296 5412 13300 5468
rect 13300 5412 13356 5468
rect 13356 5412 13360 5468
rect 13296 5408 13360 5412
rect 13376 5468 13440 5472
rect 13376 5412 13380 5468
rect 13380 5412 13436 5468
rect 13436 5412 13440 5468
rect 13376 5408 13440 5412
rect 13456 5468 13520 5472
rect 13456 5412 13460 5468
rect 13460 5412 13516 5468
rect 13516 5412 13520 5468
rect 13456 5408 13520 5412
rect 19216 5468 19280 5472
rect 19216 5412 19220 5468
rect 19220 5412 19276 5468
rect 19276 5412 19280 5468
rect 19216 5408 19280 5412
rect 19296 5468 19360 5472
rect 19296 5412 19300 5468
rect 19300 5412 19356 5468
rect 19356 5412 19360 5468
rect 19296 5408 19360 5412
rect 19376 5468 19440 5472
rect 19376 5412 19380 5468
rect 19380 5412 19436 5468
rect 19436 5412 19440 5468
rect 19376 5408 19440 5412
rect 19456 5468 19520 5472
rect 19456 5412 19460 5468
rect 19460 5412 19516 5468
rect 19516 5412 19520 5468
rect 19456 5408 19520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 10216 4924 10280 4928
rect 10216 4868 10220 4924
rect 10220 4868 10276 4924
rect 10276 4868 10280 4924
rect 10216 4864 10280 4868
rect 10296 4924 10360 4928
rect 10296 4868 10300 4924
rect 10300 4868 10356 4924
rect 10356 4868 10360 4924
rect 10296 4864 10360 4868
rect 10376 4924 10440 4928
rect 10376 4868 10380 4924
rect 10380 4868 10436 4924
rect 10436 4868 10440 4924
rect 10376 4864 10440 4868
rect 10456 4924 10520 4928
rect 10456 4868 10460 4924
rect 10460 4868 10516 4924
rect 10516 4868 10520 4924
rect 10456 4864 10520 4868
rect 16216 4924 16280 4928
rect 16216 4868 16220 4924
rect 16220 4868 16276 4924
rect 16276 4868 16280 4924
rect 16216 4864 16280 4868
rect 16296 4924 16360 4928
rect 16296 4868 16300 4924
rect 16300 4868 16356 4924
rect 16356 4868 16360 4924
rect 16296 4864 16360 4868
rect 16376 4924 16440 4928
rect 16376 4868 16380 4924
rect 16380 4868 16436 4924
rect 16436 4868 16440 4924
rect 16376 4864 16440 4868
rect 16456 4924 16520 4928
rect 16456 4868 16460 4924
rect 16460 4868 16516 4924
rect 16516 4868 16520 4924
rect 16456 4864 16520 4868
rect 7216 4380 7280 4384
rect 7216 4324 7220 4380
rect 7220 4324 7276 4380
rect 7276 4324 7280 4380
rect 7216 4320 7280 4324
rect 7296 4380 7360 4384
rect 7296 4324 7300 4380
rect 7300 4324 7356 4380
rect 7356 4324 7360 4380
rect 7296 4320 7360 4324
rect 7376 4380 7440 4384
rect 7376 4324 7380 4380
rect 7380 4324 7436 4380
rect 7436 4324 7440 4380
rect 7376 4320 7440 4324
rect 7456 4380 7520 4384
rect 7456 4324 7460 4380
rect 7460 4324 7516 4380
rect 7516 4324 7520 4380
rect 7456 4320 7520 4324
rect 13216 4380 13280 4384
rect 13216 4324 13220 4380
rect 13220 4324 13276 4380
rect 13276 4324 13280 4380
rect 13216 4320 13280 4324
rect 13296 4380 13360 4384
rect 13296 4324 13300 4380
rect 13300 4324 13356 4380
rect 13356 4324 13360 4380
rect 13296 4320 13360 4324
rect 13376 4380 13440 4384
rect 13376 4324 13380 4380
rect 13380 4324 13436 4380
rect 13436 4324 13440 4380
rect 13376 4320 13440 4324
rect 13456 4380 13520 4384
rect 13456 4324 13460 4380
rect 13460 4324 13516 4380
rect 13516 4324 13520 4380
rect 13456 4320 13520 4324
rect 19216 4380 19280 4384
rect 19216 4324 19220 4380
rect 19220 4324 19276 4380
rect 19276 4324 19280 4380
rect 19216 4320 19280 4324
rect 19296 4380 19360 4384
rect 19296 4324 19300 4380
rect 19300 4324 19356 4380
rect 19356 4324 19360 4380
rect 19296 4320 19360 4324
rect 19376 4380 19440 4384
rect 19376 4324 19380 4380
rect 19380 4324 19436 4380
rect 19436 4324 19440 4380
rect 19376 4320 19440 4324
rect 19456 4380 19520 4384
rect 19456 4324 19460 4380
rect 19460 4324 19516 4380
rect 19516 4324 19520 4380
rect 19456 4320 19520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 10216 3836 10280 3840
rect 10216 3780 10220 3836
rect 10220 3780 10276 3836
rect 10276 3780 10280 3836
rect 10216 3776 10280 3780
rect 10296 3836 10360 3840
rect 10296 3780 10300 3836
rect 10300 3780 10356 3836
rect 10356 3780 10360 3836
rect 10296 3776 10360 3780
rect 10376 3836 10440 3840
rect 10376 3780 10380 3836
rect 10380 3780 10436 3836
rect 10436 3780 10440 3836
rect 10376 3776 10440 3780
rect 10456 3836 10520 3840
rect 10456 3780 10460 3836
rect 10460 3780 10516 3836
rect 10516 3780 10520 3836
rect 10456 3776 10520 3780
rect 16216 3836 16280 3840
rect 16216 3780 16220 3836
rect 16220 3780 16276 3836
rect 16276 3780 16280 3836
rect 16216 3776 16280 3780
rect 16296 3836 16360 3840
rect 16296 3780 16300 3836
rect 16300 3780 16356 3836
rect 16356 3780 16360 3836
rect 16296 3776 16360 3780
rect 16376 3836 16440 3840
rect 16376 3780 16380 3836
rect 16380 3780 16436 3836
rect 16436 3780 16440 3836
rect 16376 3776 16440 3780
rect 16456 3836 16520 3840
rect 16456 3780 16460 3836
rect 16460 3780 16516 3836
rect 16516 3780 16520 3836
rect 16456 3776 16520 3780
rect 7216 3292 7280 3296
rect 7216 3236 7220 3292
rect 7220 3236 7276 3292
rect 7276 3236 7280 3292
rect 7216 3232 7280 3236
rect 7296 3292 7360 3296
rect 7296 3236 7300 3292
rect 7300 3236 7356 3292
rect 7356 3236 7360 3292
rect 7296 3232 7360 3236
rect 7376 3292 7440 3296
rect 7376 3236 7380 3292
rect 7380 3236 7436 3292
rect 7436 3236 7440 3292
rect 7376 3232 7440 3236
rect 7456 3292 7520 3296
rect 7456 3236 7460 3292
rect 7460 3236 7516 3292
rect 7516 3236 7520 3292
rect 7456 3232 7520 3236
rect 13216 3292 13280 3296
rect 13216 3236 13220 3292
rect 13220 3236 13276 3292
rect 13276 3236 13280 3292
rect 13216 3232 13280 3236
rect 13296 3292 13360 3296
rect 13296 3236 13300 3292
rect 13300 3236 13356 3292
rect 13356 3236 13360 3292
rect 13296 3232 13360 3236
rect 13376 3292 13440 3296
rect 13376 3236 13380 3292
rect 13380 3236 13436 3292
rect 13436 3236 13440 3292
rect 13376 3232 13440 3236
rect 13456 3292 13520 3296
rect 13456 3236 13460 3292
rect 13460 3236 13516 3292
rect 13516 3236 13520 3292
rect 13456 3232 13520 3236
rect 19216 3292 19280 3296
rect 19216 3236 19220 3292
rect 19220 3236 19276 3292
rect 19276 3236 19280 3292
rect 19216 3232 19280 3236
rect 19296 3292 19360 3296
rect 19296 3236 19300 3292
rect 19300 3236 19356 3292
rect 19356 3236 19360 3292
rect 19296 3232 19360 3236
rect 19376 3292 19440 3296
rect 19376 3236 19380 3292
rect 19380 3236 19436 3292
rect 19436 3236 19440 3292
rect 19376 3232 19440 3236
rect 19456 3292 19520 3296
rect 19456 3236 19460 3292
rect 19460 3236 19516 3292
rect 19516 3236 19520 3292
rect 19456 3232 19520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 10216 2748 10280 2752
rect 10216 2692 10220 2748
rect 10220 2692 10276 2748
rect 10276 2692 10280 2748
rect 10216 2688 10280 2692
rect 10296 2748 10360 2752
rect 10296 2692 10300 2748
rect 10300 2692 10356 2748
rect 10356 2692 10360 2748
rect 10296 2688 10360 2692
rect 10376 2748 10440 2752
rect 10376 2692 10380 2748
rect 10380 2692 10436 2748
rect 10436 2692 10440 2748
rect 10376 2688 10440 2692
rect 10456 2748 10520 2752
rect 10456 2692 10460 2748
rect 10460 2692 10516 2748
rect 10516 2692 10520 2748
rect 10456 2688 10520 2692
rect 16216 2748 16280 2752
rect 16216 2692 16220 2748
rect 16220 2692 16276 2748
rect 16276 2692 16280 2748
rect 16216 2688 16280 2692
rect 16296 2748 16360 2752
rect 16296 2692 16300 2748
rect 16300 2692 16356 2748
rect 16356 2692 16360 2748
rect 16296 2688 16360 2692
rect 16376 2748 16440 2752
rect 16376 2692 16380 2748
rect 16380 2692 16436 2748
rect 16436 2692 16440 2748
rect 16376 2688 16440 2692
rect 16456 2748 16520 2752
rect 16456 2692 16460 2748
rect 16460 2692 16516 2748
rect 16516 2692 16520 2748
rect 16456 2688 16520 2692
rect 7216 2204 7280 2208
rect 7216 2148 7220 2204
rect 7220 2148 7276 2204
rect 7276 2148 7280 2204
rect 7216 2144 7280 2148
rect 7296 2204 7360 2208
rect 7296 2148 7300 2204
rect 7300 2148 7356 2204
rect 7356 2148 7360 2204
rect 7296 2144 7360 2148
rect 7376 2204 7440 2208
rect 7376 2148 7380 2204
rect 7380 2148 7436 2204
rect 7436 2148 7440 2204
rect 7376 2144 7440 2148
rect 7456 2204 7520 2208
rect 7456 2148 7460 2204
rect 7460 2148 7516 2204
rect 7516 2148 7520 2204
rect 7456 2144 7520 2148
rect 13216 2204 13280 2208
rect 13216 2148 13220 2204
rect 13220 2148 13276 2204
rect 13276 2148 13280 2204
rect 13216 2144 13280 2148
rect 13296 2204 13360 2208
rect 13296 2148 13300 2204
rect 13300 2148 13356 2204
rect 13356 2148 13360 2204
rect 13296 2144 13360 2148
rect 13376 2204 13440 2208
rect 13376 2148 13380 2204
rect 13380 2148 13436 2204
rect 13436 2148 13440 2204
rect 13376 2144 13440 2148
rect 13456 2204 13520 2208
rect 13456 2148 13460 2204
rect 13460 2148 13516 2204
rect 13516 2148 13520 2204
rect 13456 2144 13520 2148
rect 19216 2204 19280 2208
rect 19216 2148 19220 2204
rect 19220 2148 19276 2204
rect 19276 2148 19280 2204
rect 19216 2144 19280 2148
rect 19296 2204 19360 2208
rect 19296 2148 19300 2204
rect 19300 2148 19356 2204
rect 19356 2148 19360 2204
rect 19296 2144 19360 2148
rect 19376 2204 19440 2208
rect 19376 2148 19380 2204
rect 19380 2148 19436 2204
rect 19436 2148 19440 2204
rect 19376 2144 19440 2148
rect 19456 2204 19520 2208
rect 19456 2148 19460 2204
rect 19460 2148 19516 2204
rect 19516 2148 19520 2204
rect 19456 2144 19520 2148
<< metal4 >>
rect 4208 21248 4528 21808
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 7208 21792 7528 21808
rect 7208 21728 7216 21792
rect 7280 21728 7296 21792
rect 7360 21728 7376 21792
rect 7440 21728 7456 21792
rect 7520 21728 7528 21792
rect 7208 20704 7528 21728
rect 7208 20640 7216 20704
rect 7280 20640 7296 20704
rect 7360 20640 7376 20704
rect 7440 20640 7456 20704
rect 7520 20640 7528 20704
rect 7208 19616 7528 20640
rect 7208 19552 7216 19616
rect 7280 19552 7296 19616
rect 7360 19552 7376 19616
rect 7440 19552 7456 19616
rect 7520 19552 7528 19616
rect 7208 18528 7528 19552
rect 7208 18464 7216 18528
rect 7280 18464 7296 18528
rect 7360 18464 7376 18528
rect 7440 18464 7456 18528
rect 7520 18464 7528 18528
rect 7208 17440 7528 18464
rect 7208 17376 7216 17440
rect 7280 17376 7296 17440
rect 7360 17376 7376 17440
rect 7440 17376 7456 17440
rect 7520 17376 7528 17440
rect 7208 16352 7528 17376
rect 7208 16288 7216 16352
rect 7280 16288 7296 16352
rect 7360 16288 7376 16352
rect 7440 16288 7456 16352
rect 7520 16288 7528 16352
rect 7208 15264 7528 16288
rect 7208 15200 7216 15264
rect 7280 15200 7296 15264
rect 7360 15200 7376 15264
rect 7440 15200 7456 15264
rect 7520 15200 7528 15264
rect 7208 14176 7528 15200
rect 7208 14112 7216 14176
rect 7280 14112 7296 14176
rect 7360 14112 7376 14176
rect 7440 14112 7456 14176
rect 7520 14112 7528 14176
rect 7208 13088 7528 14112
rect 7208 13024 7216 13088
rect 7280 13024 7296 13088
rect 7360 13024 7376 13088
rect 7440 13024 7456 13088
rect 7520 13024 7528 13088
rect 7208 12000 7528 13024
rect 7208 11936 7216 12000
rect 7280 11936 7296 12000
rect 7360 11936 7376 12000
rect 7440 11936 7456 12000
rect 7520 11936 7528 12000
rect 7208 10912 7528 11936
rect 7208 10848 7216 10912
rect 7280 10848 7296 10912
rect 7360 10848 7376 10912
rect 7440 10848 7456 10912
rect 7520 10848 7528 10912
rect 7208 9824 7528 10848
rect 7208 9760 7216 9824
rect 7280 9760 7296 9824
rect 7360 9760 7376 9824
rect 7440 9760 7456 9824
rect 7520 9760 7528 9824
rect 7208 8736 7528 9760
rect 7208 8672 7216 8736
rect 7280 8672 7296 8736
rect 7360 8672 7376 8736
rect 7440 8672 7456 8736
rect 7520 8672 7528 8736
rect 7208 7648 7528 8672
rect 7208 7584 7216 7648
rect 7280 7584 7296 7648
rect 7360 7584 7376 7648
rect 7440 7584 7456 7648
rect 7520 7584 7528 7648
rect 7208 6560 7528 7584
rect 7208 6496 7216 6560
rect 7280 6496 7296 6560
rect 7360 6496 7376 6560
rect 7440 6496 7456 6560
rect 7520 6496 7528 6560
rect 7208 5472 7528 6496
rect 7208 5408 7216 5472
rect 7280 5408 7296 5472
rect 7360 5408 7376 5472
rect 7440 5408 7456 5472
rect 7520 5408 7528 5472
rect 7208 4384 7528 5408
rect 7208 4320 7216 4384
rect 7280 4320 7296 4384
rect 7360 4320 7376 4384
rect 7440 4320 7456 4384
rect 7520 4320 7528 4384
rect 7208 3296 7528 4320
rect 7208 3232 7216 3296
rect 7280 3232 7296 3296
rect 7360 3232 7376 3296
rect 7440 3232 7456 3296
rect 7520 3232 7528 3296
rect 7208 2208 7528 3232
rect 7208 2144 7216 2208
rect 7280 2144 7296 2208
rect 7360 2144 7376 2208
rect 7440 2144 7456 2208
rect 7520 2144 7528 2208
rect 7208 2128 7528 2144
rect 10208 21248 10528 21808
rect 10208 21184 10216 21248
rect 10280 21184 10296 21248
rect 10360 21184 10376 21248
rect 10440 21184 10456 21248
rect 10520 21184 10528 21248
rect 10208 20160 10528 21184
rect 10208 20096 10216 20160
rect 10280 20096 10296 20160
rect 10360 20096 10376 20160
rect 10440 20096 10456 20160
rect 10520 20096 10528 20160
rect 10208 19072 10528 20096
rect 10208 19008 10216 19072
rect 10280 19008 10296 19072
rect 10360 19008 10376 19072
rect 10440 19008 10456 19072
rect 10520 19008 10528 19072
rect 10208 17984 10528 19008
rect 10208 17920 10216 17984
rect 10280 17920 10296 17984
rect 10360 17920 10376 17984
rect 10440 17920 10456 17984
rect 10520 17920 10528 17984
rect 10208 16896 10528 17920
rect 10208 16832 10216 16896
rect 10280 16832 10296 16896
rect 10360 16832 10376 16896
rect 10440 16832 10456 16896
rect 10520 16832 10528 16896
rect 10208 15808 10528 16832
rect 10208 15744 10216 15808
rect 10280 15744 10296 15808
rect 10360 15744 10376 15808
rect 10440 15744 10456 15808
rect 10520 15744 10528 15808
rect 10208 14720 10528 15744
rect 10208 14656 10216 14720
rect 10280 14656 10296 14720
rect 10360 14656 10376 14720
rect 10440 14656 10456 14720
rect 10520 14656 10528 14720
rect 10208 13632 10528 14656
rect 10208 13568 10216 13632
rect 10280 13568 10296 13632
rect 10360 13568 10376 13632
rect 10440 13568 10456 13632
rect 10520 13568 10528 13632
rect 10208 12544 10528 13568
rect 10208 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10528 12544
rect 10208 11456 10528 12480
rect 10208 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10528 11456
rect 10208 10368 10528 11392
rect 10208 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10528 10368
rect 10208 9280 10528 10304
rect 10208 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10528 9280
rect 10208 8192 10528 9216
rect 10208 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10528 8192
rect 10208 7104 10528 8128
rect 10208 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10528 7104
rect 10208 6016 10528 7040
rect 10208 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10528 6016
rect 10208 4928 10528 5952
rect 10208 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10528 4928
rect 10208 3840 10528 4864
rect 10208 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10528 3840
rect 10208 2752 10528 3776
rect 10208 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10528 2752
rect 10208 2128 10528 2688
rect 13208 21792 13528 21808
rect 13208 21728 13216 21792
rect 13280 21728 13296 21792
rect 13360 21728 13376 21792
rect 13440 21728 13456 21792
rect 13520 21728 13528 21792
rect 13208 20704 13528 21728
rect 13208 20640 13216 20704
rect 13280 20640 13296 20704
rect 13360 20640 13376 20704
rect 13440 20640 13456 20704
rect 13520 20640 13528 20704
rect 13208 19616 13528 20640
rect 13208 19552 13216 19616
rect 13280 19552 13296 19616
rect 13360 19552 13376 19616
rect 13440 19552 13456 19616
rect 13520 19552 13528 19616
rect 13208 18528 13528 19552
rect 13208 18464 13216 18528
rect 13280 18464 13296 18528
rect 13360 18464 13376 18528
rect 13440 18464 13456 18528
rect 13520 18464 13528 18528
rect 13208 17440 13528 18464
rect 13208 17376 13216 17440
rect 13280 17376 13296 17440
rect 13360 17376 13376 17440
rect 13440 17376 13456 17440
rect 13520 17376 13528 17440
rect 13208 16352 13528 17376
rect 13208 16288 13216 16352
rect 13280 16288 13296 16352
rect 13360 16288 13376 16352
rect 13440 16288 13456 16352
rect 13520 16288 13528 16352
rect 13208 15264 13528 16288
rect 13208 15200 13216 15264
rect 13280 15200 13296 15264
rect 13360 15200 13376 15264
rect 13440 15200 13456 15264
rect 13520 15200 13528 15264
rect 13208 14176 13528 15200
rect 13208 14112 13216 14176
rect 13280 14112 13296 14176
rect 13360 14112 13376 14176
rect 13440 14112 13456 14176
rect 13520 14112 13528 14176
rect 13208 13088 13528 14112
rect 13208 13024 13216 13088
rect 13280 13024 13296 13088
rect 13360 13024 13376 13088
rect 13440 13024 13456 13088
rect 13520 13024 13528 13088
rect 13208 12000 13528 13024
rect 13208 11936 13216 12000
rect 13280 11936 13296 12000
rect 13360 11936 13376 12000
rect 13440 11936 13456 12000
rect 13520 11936 13528 12000
rect 13208 10912 13528 11936
rect 13208 10848 13216 10912
rect 13280 10848 13296 10912
rect 13360 10848 13376 10912
rect 13440 10848 13456 10912
rect 13520 10848 13528 10912
rect 13208 9824 13528 10848
rect 13208 9760 13216 9824
rect 13280 9760 13296 9824
rect 13360 9760 13376 9824
rect 13440 9760 13456 9824
rect 13520 9760 13528 9824
rect 13208 8736 13528 9760
rect 13208 8672 13216 8736
rect 13280 8672 13296 8736
rect 13360 8672 13376 8736
rect 13440 8672 13456 8736
rect 13520 8672 13528 8736
rect 13208 7648 13528 8672
rect 13208 7584 13216 7648
rect 13280 7584 13296 7648
rect 13360 7584 13376 7648
rect 13440 7584 13456 7648
rect 13520 7584 13528 7648
rect 13208 6560 13528 7584
rect 13208 6496 13216 6560
rect 13280 6496 13296 6560
rect 13360 6496 13376 6560
rect 13440 6496 13456 6560
rect 13520 6496 13528 6560
rect 13208 5472 13528 6496
rect 13208 5408 13216 5472
rect 13280 5408 13296 5472
rect 13360 5408 13376 5472
rect 13440 5408 13456 5472
rect 13520 5408 13528 5472
rect 13208 4384 13528 5408
rect 13208 4320 13216 4384
rect 13280 4320 13296 4384
rect 13360 4320 13376 4384
rect 13440 4320 13456 4384
rect 13520 4320 13528 4384
rect 13208 3296 13528 4320
rect 13208 3232 13216 3296
rect 13280 3232 13296 3296
rect 13360 3232 13376 3296
rect 13440 3232 13456 3296
rect 13520 3232 13528 3296
rect 13208 2208 13528 3232
rect 13208 2144 13216 2208
rect 13280 2144 13296 2208
rect 13360 2144 13376 2208
rect 13440 2144 13456 2208
rect 13520 2144 13528 2208
rect 13208 2128 13528 2144
rect 16208 21248 16528 21808
rect 16208 21184 16216 21248
rect 16280 21184 16296 21248
rect 16360 21184 16376 21248
rect 16440 21184 16456 21248
rect 16520 21184 16528 21248
rect 16208 20160 16528 21184
rect 16208 20096 16216 20160
rect 16280 20096 16296 20160
rect 16360 20096 16376 20160
rect 16440 20096 16456 20160
rect 16520 20096 16528 20160
rect 16208 19072 16528 20096
rect 16208 19008 16216 19072
rect 16280 19008 16296 19072
rect 16360 19008 16376 19072
rect 16440 19008 16456 19072
rect 16520 19008 16528 19072
rect 16208 17984 16528 19008
rect 16208 17920 16216 17984
rect 16280 17920 16296 17984
rect 16360 17920 16376 17984
rect 16440 17920 16456 17984
rect 16520 17920 16528 17984
rect 16208 16896 16528 17920
rect 16208 16832 16216 16896
rect 16280 16832 16296 16896
rect 16360 16832 16376 16896
rect 16440 16832 16456 16896
rect 16520 16832 16528 16896
rect 16208 15808 16528 16832
rect 16208 15744 16216 15808
rect 16280 15744 16296 15808
rect 16360 15744 16376 15808
rect 16440 15744 16456 15808
rect 16520 15744 16528 15808
rect 16208 14720 16528 15744
rect 16208 14656 16216 14720
rect 16280 14656 16296 14720
rect 16360 14656 16376 14720
rect 16440 14656 16456 14720
rect 16520 14656 16528 14720
rect 16208 13632 16528 14656
rect 16208 13568 16216 13632
rect 16280 13568 16296 13632
rect 16360 13568 16376 13632
rect 16440 13568 16456 13632
rect 16520 13568 16528 13632
rect 16208 12544 16528 13568
rect 16208 12480 16216 12544
rect 16280 12480 16296 12544
rect 16360 12480 16376 12544
rect 16440 12480 16456 12544
rect 16520 12480 16528 12544
rect 16208 11456 16528 12480
rect 16208 11392 16216 11456
rect 16280 11392 16296 11456
rect 16360 11392 16376 11456
rect 16440 11392 16456 11456
rect 16520 11392 16528 11456
rect 16208 10368 16528 11392
rect 16208 10304 16216 10368
rect 16280 10304 16296 10368
rect 16360 10304 16376 10368
rect 16440 10304 16456 10368
rect 16520 10304 16528 10368
rect 16208 9280 16528 10304
rect 16208 9216 16216 9280
rect 16280 9216 16296 9280
rect 16360 9216 16376 9280
rect 16440 9216 16456 9280
rect 16520 9216 16528 9280
rect 16208 8192 16528 9216
rect 16208 8128 16216 8192
rect 16280 8128 16296 8192
rect 16360 8128 16376 8192
rect 16440 8128 16456 8192
rect 16520 8128 16528 8192
rect 16208 7104 16528 8128
rect 16208 7040 16216 7104
rect 16280 7040 16296 7104
rect 16360 7040 16376 7104
rect 16440 7040 16456 7104
rect 16520 7040 16528 7104
rect 16208 6016 16528 7040
rect 16208 5952 16216 6016
rect 16280 5952 16296 6016
rect 16360 5952 16376 6016
rect 16440 5952 16456 6016
rect 16520 5952 16528 6016
rect 16208 4928 16528 5952
rect 16208 4864 16216 4928
rect 16280 4864 16296 4928
rect 16360 4864 16376 4928
rect 16440 4864 16456 4928
rect 16520 4864 16528 4928
rect 16208 3840 16528 4864
rect 16208 3776 16216 3840
rect 16280 3776 16296 3840
rect 16360 3776 16376 3840
rect 16440 3776 16456 3840
rect 16520 3776 16528 3840
rect 16208 2752 16528 3776
rect 16208 2688 16216 2752
rect 16280 2688 16296 2752
rect 16360 2688 16376 2752
rect 16440 2688 16456 2752
rect 16520 2688 16528 2752
rect 16208 2128 16528 2688
rect 19208 21792 19528 21808
rect 19208 21728 19216 21792
rect 19280 21728 19296 21792
rect 19360 21728 19376 21792
rect 19440 21728 19456 21792
rect 19520 21728 19528 21792
rect 19208 20704 19528 21728
rect 19208 20640 19216 20704
rect 19280 20640 19296 20704
rect 19360 20640 19376 20704
rect 19440 20640 19456 20704
rect 19520 20640 19528 20704
rect 19208 19616 19528 20640
rect 19208 19552 19216 19616
rect 19280 19552 19296 19616
rect 19360 19552 19376 19616
rect 19440 19552 19456 19616
rect 19520 19552 19528 19616
rect 19208 18528 19528 19552
rect 19208 18464 19216 18528
rect 19280 18464 19296 18528
rect 19360 18464 19376 18528
rect 19440 18464 19456 18528
rect 19520 18464 19528 18528
rect 19208 17440 19528 18464
rect 19208 17376 19216 17440
rect 19280 17376 19296 17440
rect 19360 17376 19376 17440
rect 19440 17376 19456 17440
rect 19520 17376 19528 17440
rect 19208 16352 19528 17376
rect 19208 16288 19216 16352
rect 19280 16288 19296 16352
rect 19360 16288 19376 16352
rect 19440 16288 19456 16352
rect 19520 16288 19528 16352
rect 19208 15264 19528 16288
rect 19208 15200 19216 15264
rect 19280 15200 19296 15264
rect 19360 15200 19376 15264
rect 19440 15200 19456 15264
rect 19520 15200 19528 15264
rect 19208 14176 19528 15200
rect 19208 14112 19216 14176
rect 19280 14112 19296 14176
rect 19360 14112 19376 14176
rect 19440 14112 19456 14176
rect 19520 14112 19528 14176
rect 19208 13088 19528 14112
rect 19208 13024 19216 13088
rect 19280 13024 19296 13088
rect 19360 13024 19376 13088
rect 19440 13024 19456 13088
rect 19520 13024 19528 13088
rect 19208 12000 19528 13024
rect 19208 11936 19216 12000
rect 19280 11936 19296 12000
rect 19360 11936 19376 12000
rect 19440 11936 19456 12000
rect 19520 11936 19528 12000
rect 19208 10912 19528 11936
rect 19208 10848 19216 10912
rect 19280 10848 19296 10912
rect 19360 10848 19376 10912
rect 19440 10848 19456 10912
rect 19520 10848 19528 10912
rect 19208 9824 19528 10848
rect 19208 9760 19216 9824
rect 19280 9760 19296 9824
rect 19360 9760 19376 9824
rect 19440 9760 19456 9824
rect 19520 9760 19528 9824
rect 19208 8736 19528 9760
rect 19208 8672 19216 8736
rect 19280 8672 19296 8736
rect 19360 8672 19376 8736
rect 19440 8672 19456 8736
rect 19520 8672 19528 8736
rect 19208 7648 19528 8672
rect 19208 7584 19216 7648
rect 19280 7584 19296 7648
rect 19360 7584 19376 7648
rect 19440 7584 19456 7648
rect 19520 7584 19528 7648
rect 19208 6560 19528 7584
rect 19208 6496 19216 6560
rect 19280 6496 19296 6560
rect 19360 6496 19376 6560
rect 19440 6496 19456 6560
rect 19520 6496 19528 6560
rect 19208 5472 19528 6496
rect 19208 5408 19216 5472
rect 19280 5408 19296 5472
rect 19360 5408 19376 5472
rect 19440 5408 19456 5472
rect 19520 5408 19528 5472
rect 19208 4384 19528 5408
rect 19208 4320 19216 4384
rect 19280 4320 19296 4384
rect 19360 4320 19376 4384
rect 19440 4320 19456 4384
rect 19520 4320 19528 4384
rect 19208 3296 19528 4320
rect 19208 3232 19216 3296
rect 19280 3232 19296 3296
rect 19360 3232 19376 3296
rect 19440 3232 19456 3296
rect 19520 3232 19528 3296
rect 19208 2208 19528 3232
rect 19208 2144 19216 2208
rect 19280 2144 19296 2208
rect 19360 2144 19376 2208
rect 19440 2144 19456 2208
rect 19520 2144 19528 2208
rect 19208 2128 19528 2144
use sky130_fd_sc_hd__and4_1  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 17296 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 15456 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _169_
timestamp 1692646696
transform 1 0 14076 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _170_
timestamp 1692646696
transform -1 0 16192 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1692646696
transform 1 0 15824 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 19044 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 15916 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _174_
timestamp 1692646696
transform 1 0 13800 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _175_
timestamp 1692646696
transform 1 0 15824 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _176_
timestamp 1692646696
transform 1 0 16284 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 18032 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 17204 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _179_
timestamp 1692646696
transform 1 0 14536 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _180_
timestamp 1692646696
transform -1 0 14536 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _181_
timestamp 1692646696
transform 1 0 12052 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _182_
timestamp 1692646696
transform 1 0 14076 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _183_
timestamp 1692646696
transform 1 0 14168 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _184_
timestamp 1692646696
transform 1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _185_
timestamp 1692646696
transform 1 0 14628 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _186_
timestamp 1692646696
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _187_
timestamp 1692646696
transform 1 0 15456 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _188_
timestamp 1692646696
transform 1 0 14628 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _189_
timestamp 1692646696
transform 1 0 15640 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _190_
timestamp 1692646696
transform -1 0 16008 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _191_
timestamp 1692646696
transform 1 0 18492 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _192_
timestamp 1692646696
transform 1 0 16100 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _193_
timestamp 1692646696
transform 1 0 16928 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _194_
timestamp 1692646696
transform -1 0 19872 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _195_
timestamp 1692646696
transform 1 0 17204 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _196_
timestamp 1692646696
transform -1 0 18492 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _197_
timestamp 1692646696
transform 1 0 16652 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _198_
timestamp 1692646696
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _199_
timestamp 1692646696
transform 1 0 19872 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _200_
timestamp 1692646696
transform -1 0 17848 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _201_
timestamp 1692646696
transform 1 0 17388 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _202_
timestamp 1692646696
transform 1 0 18124 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _203_
timestamp 1692646696
transform 1 0 19228 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _204_
timestamp 1692646696
transform 1 0 16100 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _205_
timestamp 1692646696
transform -1 0 18308 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _206_
timestamp 1692646696
transform -1 0 19872 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _207_
timestamp 1692646696
transform 1 0 17848 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _208_
timestamp 1692646696
transform -1 0 19136 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _209_
timestamp 1692646696
transform 1 0 16928 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _210_
timestamp 1692646696
transform 1 0 17756 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _211_
timestamp 1692646696
transform -1 0 19780 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _212_
timestamp 1692646696
transform -1 0 18584 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _213_
timestamp 1692646696
transform -1 0 17664 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _214_
timestamp 1692646696
transform 1 0 17664 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _216_
timestamp 1692646696
transform 1 0 16928 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 17572 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _218_
timestamp 1692646696
transform 1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 9660 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 13064 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1692646696
transform 1 0 13616 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 4048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1692646696
transform 1 0 6440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _224_
timestamp 1692646696
transform 1 0 3772 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1692646696
transform 1 0 6624 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _226_
timestamp 1692646696
transform -1 0 7360 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _227_
timestamp 1692646696
transform 1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1692646696
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _229_
timestamp 1692646696
transform 1 0 4416 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1692646696
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _232_
timestamp 1692646696
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _233_
timestamp 1692646696
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1692646696
transform -1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _235_
timestamp 1692646696
transform -1 0 12236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _236_
timestamp 1692646696
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _237_
timestamp 1692646696
transform -1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 10396 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 11040 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1692646696
transform -1 0 11960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _241_
timestamp 1692646696
transform -1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _242_
timestamp 1692646696
transform 1 0 12328 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1692646696
transform 1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _244_
timestamp 1692646696
transform 1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _245_
timestamp 1692646696
transform 1 0 11960 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1692646696
transform -1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _247_
timestamp 1692646696
transform -1 0 3312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1692646696
transform 1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp 1692646696
transform 1 0 3496 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _250_
timestamp 1692646696
transform 1 0 1656 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1692646696
transform 1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _252_
timestamp 1692646696
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _253_
timestamp 1692646696
transform 1 0 3864 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1692646696
transform 1 0 4692 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _255_
timestamp 1692646696
transform 1 0 1472 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _256_
timestamp 1692646696
transform -1 0 7452 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1692646696
transform -1 0 6716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _258_
timestamp 1692646696
transform 1 0 7452 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1692646696
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _260_
timestamp 1692646696
transform -1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _261_
timestamp 1692646696
transform -1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _262_
timestamp 1692646696
transform 1 0 10764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1692646696
transform -1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _264_
timestamp 1692646696
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _265_
timestamp 1692646696
transform 1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 7360 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _267_
timestamp 1692646696
transform -1 0 9936 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 9476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _269_
timestamp 1692646696
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _270_
timestamp 1692646696
transform 1 0 9936 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _271_
timestamp 1692646696
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _272_
timestamp 1692646696
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 10580 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 10396 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 9936 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1692646696
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 10396 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _278_
timestamp 1692646696
transform 1 0 11500 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 11408 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _280_
timestamp 1692646696
transform -1 0 12696 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _281_
timestamp 1692646696
transform -1 0 11408 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _282_
timestamp 1692646696
transform 1 0 10764 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 10488 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 10212 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _285_
timestamp 1692646696
transform -1 0 10120 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1692646696
transform -1 0 11684 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _287_
timestamp 1692646696
transform -1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1692646696
transform -1 0 11960 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _289_
timestamp 1692646696
transform -1 0 11960 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1692646696
transform -1 0 10028 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _291_
timestamp 1692646696
transform -1 0 11224 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _292_
timestamp 1692646696
transform 1 0 1380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _293_
timestamp 1692646696
transform 1 0 3772 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _294_
timestamp 1692646696
transform -1 0 4600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _295_
timestamp 1692646696
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _296_
timestamp 1692646696
transform 1 0 4784 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _297_
timestamp 1692646696
transform 1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _298_
timestamp 1692646696
transform -1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _299_
timestamp 1692646696
transform -1 0 5152 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _300_
timestamp 1692646696
transform 1 0 6072 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _301_
timestamp 1692646696
transform -1 0 6256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1692646696
transform 1 0 6256 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1692646696
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _304_
timestamp 1692646696
transform 1 0 6900 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _305_
timestamp 1692646696
transform 1 0 6900 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1692646696
transform -1 0 7636 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _307_
timestamp 1692646696
transform 1 0 7912 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1692646696
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1692646696
transform -1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _310_
timestamp 1692646696
transform -1 0 6164 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _311_
timestamp 1692646696
transform 1 0 3956 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _312_
timestamp 1692646696
transform 1 0 5612 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _314_
timestamp 1692646696
transform -1 0 8832 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1692646696
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _316_
timestamp 1692646696
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _317_
timestamp 1692646696
transform 1 0 8740 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1692646696
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1692646696
transform 1 0 12788 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1692646696
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1692646696
transform 1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _322_
timestamp 1692646696
transform 1 0 9752 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1692646696
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1692646696
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325_
timestamp 1692646696
transform -1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1692646696
transform -1 0 2300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1692646696
transform 1 0 1748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1692646696
transform 1 0 4416 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _329_
timestamp 1692646696
transform -1 0 9752 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _331_
timestamp 1692646696
transform 1 0 6716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1692646696
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _334_
timestamp 1692646696
transform 1 0 4876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 4140 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 9660 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _337_
timestamp 1692646696
transform 1 0 4692 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _338_
timestamp 1692646696
transform 1 0 5152 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 6256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 5152 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _341_
timestamp 1692646696
transform -1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _342_
timestamp 1692646696
transform 1 0 6348 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 4508 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _345_
timestamp 1692646696
transform 1 0 3864 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _346_
timestamp 1692646696
transform 1 0 4968 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 5980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _348_
timestamp 1692646696
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _349_
timestamp 1692646696
transform -1 0 5152 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _350_
timestamp 1692646696
transform 1 0 6256 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _351_
timestamp 1692646696
transform 1 0 5612 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _352_
timestamp 1692646696
transform 1 0 6900 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _353_
timestamp 1692646696
transform 1 0 7360 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1692646696
transform -1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _355_
timestamp 1692646696
transform -1 0 7360 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _356_
timestamp 1692646696
transform -1 0 8832 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 7912 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1692646696
transform 1 0 8648 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359_
timestamp 1692646696
transform 1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _360_
timestamp 1692646696
transform 1 0 3772 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  _361_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 7636 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 6164 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _363_
timestamp 1692646696
transform 1 0 7728 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _364_
timestamp 1692646696
transform -1 0 10764 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _365_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 8280 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _366_
timestamp 1692646696
transform 1 0 8004 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _367_
timestamp 1692646696
transform 1 0 8740 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _368_
timestamp 1692646696
transform 1 0 10580 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _369_
timestamp 1692646696
transform 1 0 8556 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _370_
timestamp 1692646696
transform 1 0 11132 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _371_
timestamp 1692646696
transform 1 0 11408 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _372_
timestamp 1692646696
transform 1 0 11500 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _373_
timestamp 1692646696
transform -1 0 11960 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _374_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 11960 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _375_
timestamp 1692646696
transform 1 0 9936 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _376_
timestamp 1692646696
transform 1 0 10028 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _377_
timestamp 1692646696
transform 1 0 13800 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _378_
timestamp 1692646696
transform 1 0 11960 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _379_
timestamp 1692646696
transform 1 0 11776 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _380_
timestamp 1692646696
transform 1 0 10580 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1692646696
transform 1 0 14168 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1692646696
transform 1 0 12328 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1692646696
transform 1 0 14720 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1692646696
transform 1 0 12880 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _385_
timestamp 1692646696
transform 1 0 14168 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _386_
timestamp 1692646696
transform 1 0 12328 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _387_
timestamp 1692646696
transform 1 0 10120 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _388_
timestamp 1692646696
transform -1 0 10764 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1692646696
transform 1 0 3496 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1692646696
transform 1 0 4232 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _391_
timestamp 1692646696
transform 1 0 1840 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _392_
timestamp 1692646696
transform 1 0 3772 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _393__22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 4692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1692646696
transform 1 0 3864 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1692646696
transform 1 0 5796 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1692646696
transform 1 0 6808 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1692646696
transform 1 0 2576 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1692646696
transform 1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1692646696
transform 1 0 1380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1692646696
transform 1 0 1840 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1692646696
transform 1 0 1380 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1692646696
transform 1 0 2024 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1692646696
transform 1 0 3772 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1692646696
transform -1 0 6256 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _404_
timestamp 1692646696
transform 1 0 1840 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _405_
timestamp 1692646696
transform 1 0 2300 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _406_
timestamp 1692646696
transform 1 0 4416 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _407_
timestamp 1692646696
transform -1 0 8096 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _408_
timestamp 1692646696
transform 1 0 1840 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _409_
timestamp 1692646696
transform 1 0 3772 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _410_
timestamp 1692646696
transform 1 0 6348 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _411_
timestamp 1692646696
transform 1 0 6440 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _412_
timestamp 1692646696
transform 1 0 8556 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _413_
timestamp 1692646696
transform 1 0 4784 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _414_
timestamp 1692646696
transform 1 0 6624 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _415_
timestamp 1692646696
transform 1 0 6348 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _416_
timestamp 1692646696
transform 1 0 6716 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 1656 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _418_
timestamp 1692646696
transform 1 0 1840 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _419_
timestamp 1692646696
transform 1 0 3220 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _420_
timestamp 1692646696
transform 1 0 5704 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _421_
timestamp 1692646696
transform 1 0 4324 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _422_
timestamp 1692646696
transform -1 0 7912 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _423_
timestamp 1692646696
transform -1 0 7912 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _424_
timestamp 1692646696
transform 1 0 8924 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _425_
timestamp 1692646696
transform 1 0 16928 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _426_
timestamp 1692646696
transform -1 0 19136 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _427_
timestamp 1692646696
transform -1 0 20332 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _428_
timestamp 1692646696
transform 1 0 17940 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _429_
timestamp 1692646696
transform 1 0 16652 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _430_
timestamp 1692646696
transform 1 0 15640 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _431_
timestamp 1692646696
transform 1 0 14904 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _432_
timestamp 1692646696
transform -1 0 15824 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _433_
timestamp 1692646696
transform 1 0 14076 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _434_
timestamp 1692646696
transform 1 0 13340 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _435_
timestamp 1692646696
transform 1 0 12420 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _436_
timestamp 1692646696
transform -1 0 13984 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _437_
timestamp 1692646696
transform -1 0 14904 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _438_
timestamp 1692646696
transform -1 0 16744 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _439_
timestamp 1692646696
transform 1 0 14904 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _440_
timestamp 1692646696
transform 1 0 14076 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _441_
timestamp 1692646696
transform 1 0 14996 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _442_
timestamp 1692646696
transform -1 0 15824 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _443_
timestamp 1692646696
transform 1 0 14076 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _444_
timestamp 1692646696
transform 1 0 12880 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _445_
timestamp 1692646696
transform -1 0 14260 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _446_
timestamp 1692646696
transform -1 0 15456 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _447_
timestamp 1692646696
transform -1 0 15640 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _448_
timestamp 1692646696
transform 1 0 12328 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _449_
timestamp 1692646696
transform 1 0 11408 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _450_
timestamp 1692646696
transform -1 0 13064 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _451_
timestamp 1692646696
transform 1 0 10488 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _452_
timestamp 1692646696
transform -1 0 12236 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _453_
timestamp 1692646696
transform -1 0 13064 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _454_
timestamp 1692646696
transform -1 0 15640 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _455_
timestamp 1692646696
transform 1 0 13064 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _456_
timestamp 1692646696
transform -1 0 13984 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _457_
timestamp 1692646696
transform 1 0 16560 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _458_
timestamp 1692646696
transform -1 0 20148 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _459_
timestamp 1692646696
transform 1 0 17020 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _460_
timestamp 1692646696
transform -1 0 20056 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _461_
timestamp 1692646696
transform 1 0 17848 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _462_
timestamp 1692646696
transform -1 0 19136 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _463_
timestamp 1692646696
transform -1 0 20056 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _464_
timestamp 1692646696
transform -1 0 19688 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _465_
timestamp 1692646696
transform 1 0 18216 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _466_
timestamp 1692646696
transform -1 0 18216 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _467_
timestamp 1692646696
transform 1 0 16652 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _468_
timestamp 1692646696
transform 1 0 15364 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _469_
timestamp 1692646696
transform 1 0 14904 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _470_
timestamp 1692646696
transform -1 0 17204 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _471_
timestamp 1692646696
transform 1 0 14720 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _472_
timestamp 1692646696
transform 1 0 14076 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _473_
timestamp 1692646696
transform -1 0 18400 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _474_
timestamp 1692646696
transform -1 0 19964 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _475_
timestamp 1692646696
transform -1 0 20240 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _476_
timestamp 1692646696
transform -1 0 20424 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _477_
timestamp 1692646696
transform 1 0 17572 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _478_
timestamp 1692646696
transform -1 0 19780 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _479_
timestamp 1692646696
transform 1 0 18216 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _480_
timestamp 1692646696
transform -1 0 20516 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _481_
timestamp 1692646696
transform 1 0 18216 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _482_
timestamp 1692646696
transform -1 0 19136 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _483_
timestamp 1692646696
transform 1 0 17296 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _484_
timestamp 1692646696
transform 1 0 16652 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _485_
timestamp 1692646696
transform 1 0 15548 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _486_
timestamp 1692646696
transform -1 0 17296 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _487_
timestamp 1692646696
transform -1 0 18216 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _488_
timestamp 1692646696
transform 1 0 15364 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1692646696
transform 1 0 7728 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1692646696
transform 1 0 8924 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 1692646696
transform 1 0 9568 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 1692646696
transform 1 0 11500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 1692646696
transform 1 0 6900 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1692646696
transform 1 0 7912 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1692646696
transform 1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 1692646696
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__A
timestamp 1692646696
transform 1 0 8740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__A
timestamp 1692646696
transform 1 0 4416 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__CLK
timestamp 1692646696
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__CLK
timestamp 1692646696
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__CLK
timestamp 1692646696
transform 1 0 7544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__CLK
timestamp 1692646696
transform 1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__CLK
timestamp 1692646696
transform 1 0 8096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__CLK
timestamp 1692646696
transform 1 0 7820 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__CLK
timestamp 1692646696
transform 1 0 8556 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__CLK
timestamp 1692646696
transform 1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__CLK
timestamp 1692646696
transform 1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__CLK
timestamp 1692646696
transform 1 0 10948 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__CLK
timestamp 1692646696
transform 1 0 10948 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__CLK
timestamp 1692646696
transform -1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__CLK
timestamp 1692646696
transform 1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__CLK
timestamp 1692646696
transform 1 0 2392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__CLK
timestamp 1692646696
transform 1 0 3680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__CLK
timestamp 1692646696
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__CLK
timestamp 1692646696
transform 1 0 4232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__CLK
timestamp 1692646696
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__CLK
timestamp 1692646696
transform 1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__CLK
timestamp 1692646696
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__CLK
timestamp 1692646696
transform 1 0 6164 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__CLK
timestamp 1692646696
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__CLK
timestamp 1692646696
transform 1 0 7728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__CLK
timestamp 1692646696
transform 1 0 3220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__CLK
timestamp 1692646696
transform 1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__CLK
timestamp 1692646696
transform 1 0 2852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__CLK
timestamp 1692646696
transform 1 0 5520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__CLK
timestamp 1692646696
transform 1 0 4140 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__CLK
timestamp 1692646696
transform 1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__CLK
timestamp 1692646696
transform 1 0 5796 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__CLK
timestamp 1692646696
transform -1 0 8832 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__CLK
timestamp 1692646696
transform 1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__CLK
timestamp 1692646696
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__CLK
timestamp 1692646696
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__CLK
timestamp 1692646696
transform 1 0 17112 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__CLK
timestamp 1692646696
transform 1 0 16652 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__CLK
timestamp 1692646696
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__CLK
timestamp 1692646696
transform 1 0 14720 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__CLK
timestamp 1692646696
transform 1 0 14076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__CLK
timestamp 1692646696
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__CLK
timestamp 1692646696
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__CLK
timestamp 1692646696
transform 1 0 12236 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__CLK
timestamp 1692646696
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__CLK
timestamp 1692646696
transform 1 0 13156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__CLK
timestamp 1692646696
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__CLK
timestamp 1692646696
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__CLK
timestamp 1692646696
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__CLK
timestamp 1692646696
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__CLK
timestamp 1692646696
transform 1 0 14076 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__CLK
timestamp 1692646696
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__CLK
timestamp 1692646696
transform 1 0 12696 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__CLK
timestamp 1692646696
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__CLK
timestamp 1692646696
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__CLK
timestamp 1692646696
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__CLK
timestamp 1692646696
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__CLK
timestamp 1692646696
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__CLK
timestamp 1692646696
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__CLK
timestamp 1692646696
transform 1 0 10304 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__CLK
timestamp 1692646696
transform 1 0 10488 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__CLK
timestamp 1692646696
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__CLK
timestamp 1692646696
transform 1 0 13800 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__CLK
timestamp 1692646696
transform 1 0 12880 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__CLK
timestamp 1692646696
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__CLK
timestamp 1692646696
transform 1 0 16376 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__CLK
timestamp 1692646696
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__CLK
timestamp 1692646696
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__CLK
timestamp 1692646696
transform 1 0 18308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__CLK
timestamp 1692646696
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__CLK
timestamp 1692646696
transform 1 0 17020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__CLK
timestamp 1692646696
transform 1 0 18308 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__CLK
timestamp 1692646696
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__CLK
timestamp 1692646696
transform 1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__CLK
timestamp 1692646696
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__CLK
timestamp 1692646696
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__CLK
timestamp 1692646696
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__CLK
timestamp 1692646696
transform 1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__CLK
timestamp 1692646696
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__471__CLK
timestamp 1692646696
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__472__CLK
timestamp 1692646696
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__473__CLK
timestamp 1692646696
transform 1 0 16652 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__474__CLK
timestamp 1692646696
transform 1 0 18216 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__475__CLK
timestamp 1692646696
transform 1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__476__CLK
timestamp 1692646696
transform 1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__477__CLK
timestamp 1692646696
transform 1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__478__CLK
timestamp 1692646696
transform 1 0 18032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__479__CLK
timestamp 1692646696
transform 1 0 18492 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__480__CLK
timestamp 1692646696
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__481__CLK
timestamp 1692646696
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__482__CLK
timestamp 1692646696
transform 1 0 17388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__483__CLK
timestamp 1692646696
transform 1 0 17112 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__484__CLK
timestamp 1692646696
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__485__CLK
timestamp 1692646696
transform 1 0 15364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__486__CLK
timestamp 1692646696
transform 1 0 15548 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__487__CLK
timestamp 1692646696
transform 1 0 16836 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__488__CLK
timestamp 1692646696
transform 1 0 15180 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_4  fanout14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 1692646696
transform -1 0 6808 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 1692646696
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout17
timestamp 1692646696
transform -1 0 8832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout18
timestamp 1692646696
transform -1 0 10304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1692646696
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1692646696
transform 1 0 9936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout21
timestamp 1692646696
transform -1 0 13524 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1692646696
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1692646696
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1692646696
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1692646696
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1692646696
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97
timestamp 1692646696
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1692646696
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1692646696
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_121 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_126
timestamp 1692646696
transform 1 0 12696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_130
timestamp 1692646696
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1692646696
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1692646696
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153
timestamp 1692646696
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_161 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1692646696
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1692646696
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1692646696
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1692646696
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1692646696
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_209
timestamp 1692646696
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1692646696
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_15
timestamp 1692646696
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_23
timestamp 1692646696
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_46
timestamp 1692646696
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1692646696
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1692646696
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_69
timestamp 1692646696
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_75
timestamp 1692646696
transform 1 0 8004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_83
timestamp 1692646696
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1692646696
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1692646696
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_121
timestamp 1692646696
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_162
timestamp 1692646696
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1692646696
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1692646696
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1692646696
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_205
timestamp 1692646696
transform 1 0 19964 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1692646696
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1692646696
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1692646696
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1692646696
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_54
timestamp 1692646696
transform 1 0 6072 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_62
timestamp 1692646696
transform 1 0 6808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1692646696
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_93
timestamp 1692646696
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_97
timestamp 1692646696
transform 1 0 10028 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_134
timestamp 1692646696
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1692646696
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1692646696
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1692646696
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1692646696
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1692646696
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1692646696
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1692646696
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_209
timestamp 1692646696
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1692646696
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1692646696
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1692646696
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1692646696
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1692646696
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1692646696
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1692646696
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_69
timestamp 1692646696
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1692646696
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1692646696
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_116
timestamp 1692646696
transform 1 0 11776 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_127
timestamp 1692646696
transform 1 0 12788 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_139
timestamp 1692646696
transform 1 0 13892 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_151
timestamp 1692646696
transform 1 0 14996 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_163
timestamp 1692646696
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1692646696
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1692646696
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1692646696
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1692646696
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_205
timestamp 1692646696
transform 1 0 19964 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1692646696
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1692646696
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1692646696
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_29
timestamp 1692646696
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_35
timestamp 1692646696
transform 1 0 4324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_43
timestamp 1692646696
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_51
timestamp 1692646696
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_58
timestamp 1692646696
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_70
timestamp 1692646696
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1692646696
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_93
timestamp 1692646696
transform 1 0 9660 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_105
timestamp 1692646696
transform 1 0 10764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_117
timestamp 1692646696
transform 1 0 11868 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_125
timestamp 1692646696
transform 1 0 12604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_131
timestamp 1692646696
transform 1 0 13156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1692646696
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_145
timestamp 1692646696
transform 1 0 14444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_157
timestamp 1692646696
transform 1 0 15548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_169
timestamp 1692646696
transform 1 0 16652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1692646696
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1692646696
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1692646696
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_209
timestamp 1692646696
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1692646696
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_15
timestamp 1692646696
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_24
timestamp 1692646696
transform 1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_77
timestamp 1692646696
transform 1 0 8188 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_94
timestamp 1692646696
transform 1 0 9752 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_118
timestamp 1692646696
transform 1 0 11960 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1692646696
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_181
timestamp 1692646696
transform 1 0 17756 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_202
timestamp 1692646696
transform 1 0 19688 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_6
timestamp 1692646696
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_49
timestamp 1692646696
transform 1 0 5612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_78
timestamp 1692646696
transform 1 0 8280 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1692646696
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 1692646696
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_93
timestamp 1692646696
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_121
timestamp 1692646696
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1692646696
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1692646696
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1692646696
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1692646696
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_165
timestamp 1692646696
transform 1 0 16284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_186
timestamp 1692646696
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1692646696
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1692646696
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_209
timestamp 1692646696
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1692646696
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_15
timestamp 1692646696
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_19
timestamp 1692646696
transform 1 0 2852 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_24
timestamp 1692646696
transform 1 0 3312 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_36
timestamp 1692646696
transform 1 0 4416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_48
timestamp 1692646696
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1692646696
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_69
timestamp 1692646696
transform 1 0 7452 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_92
timestamp 1692646696
transform 1 0 9568 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_100
timestamp 1692646696
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1692646696
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_113
timestamp 1692646696
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_121
timestamp 1692646696
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_162
timestamp 1692646696
transform 1 0 16008 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_203
timestamp 1692646696
transform 1 0 19780 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1692646696
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1692646696
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1692646696
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1692646696
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1692646696
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_53
timestamp 1692646696
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_57
timestamp 1692646696
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 1692646696
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1692646696
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1692646696
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1692646696
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1692646696
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_121
timestamp 1692646696
transform 1 0 12236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_130
timestamp 1692646696
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1692646696
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1692646696
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_185
timestamp 1692646696
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1692646696
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1692646696
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1692646696
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_209
timestamp 1692646696
transform 1 0 20332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1692646696
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1692646696
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_27
timestamp 1692646696
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_30
timestamp 1692646696
transform 1 0 3864 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_36
timestamp 1692646696
transform 1 0 4416 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1692646696
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_77
timestamp 1692646696
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_93
timestamp 1692646696
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_100
timestamp 1692646696
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_116
timestamp 1692646696
transform 1 0 11776 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_128
timestamp 1692646696
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_140
timestamp 1692646696
transform 1 0 13984 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1692646696
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1692646696
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_181
timestamp 1692646696
transform 1 0 17756 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_206
timestamp 1692646696
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_210
timestamp 1692646696
transform 1 0 20424 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1692646696
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_7
timestamp 1692646696
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_59
timestamp 1692646696
transform 1 0 6532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_73
timestamp 1692646696
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_105
timestamp 1692646696
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_114
timestamp 1692646696
transform 1 0 11592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1692646696
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 1692646696
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_145
timestamp 1692646696
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_165
timestamp 1692646696
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_175
timestamp 1692646696
transform 1 0 17204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_210
timestamp 1692646696
transform 1 0 20424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_16
timestamp 1692646696
transform 1 0 2576 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_24
timestamp 1692646696
transform 1 0 3312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_29
timestamp 1692646696
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1692646696
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1692646696
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_78
timestamp 1692646696
transform 1 0 8280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_94
timestamp 1692646696
transform 1 0 9752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_100
timestamp 1692646696
transform 1 0 10304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1692646696
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_158
timestamp 1692646696
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_162
timestamp 1692646696
transform 1 0 16008 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_174
timestamp 1692646696
transform 1 0 17112 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_180
timestamp 1692646696
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_199
timestamp 1692646696
transform 1 0 19412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_3
timestamp 1692646696
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_14
timestamp 1692646696
transform 1 0 2392 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1692646696
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1692646696
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_43
timestamp 1692646696
transform 1 0 5060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_55
timestamp 1692646696
transform 1 0 6164 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_58
timestamp 1692646696
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_62
timestamp 1692646696
transform 1 0 6808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_69
timestamp 1692646696
transform 1 0 7452 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_74
timestamp 1692646696
transform 1 0 7912 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1692646696
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_97
timestamp 1692646696
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_123
timestamp 1692646696
transform 1 0 12420 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_135
timestamp 1692646696
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_175
timestamp 1692646696
transform 1 0 17204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_182
timestamp 1692646696
transform 1 0 17848 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_186
timestamp 1692646696
transform 1 0 18216 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1692646696
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_209
timestamp 1692646696
transform 1 0 20332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1692646696
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_13
timestamp 1692646696
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_17
timestamp 1692646696
transform 1 0 2668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_25
timestamp 1692646696
transform 1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_30
timestamp 1692646696
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_42
timestamp 1692646696
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_60
timestamp 1692646696
transform 1 0 6624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_64
timestamp 1692646696
transform 1 0 6992 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_101
timestamp 1692646696
transform 1 0 10396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1692646696
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1692646696
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1692646696
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1692646696
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_149
timestamp 1692646696
transform 1 0 14812 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_155
timestamp 1692646696
transform 1 0 15364 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_158
timestamp 1692646696
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1692646696
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_169
timestamp 1692646696
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_182
timestamp 1692646696
transform 1 0 17848 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_206
timestamp 1692646696
transform 1 0 20056 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_210
timestamp 1692646696
transform 1 0 20424 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1692646696
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_38
timestamp 1692646696
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_55
timestamp 1692646696
transform 1 0 6164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_76
timestamp 1692646696
transform 1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_94
timestamp 1692646696
transform 1 0 9752 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_118
timestamp 1692646696
transform 1 0 11960 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_130
timestamp 1692646696
transform 1 0 13064 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_133
timestamp 1692646696
transform 1 0 13340 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_137
timestamp 1692646696
transform 1 0 13708 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_158
timestamp 1692646696
transform 1 0 15640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1692646696
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1692646696
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1692646696
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_64
timestamp 1692646696
transform 1 0 6992 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_68
timestamp 1692646696
transform 1 0 7360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_92
timestamp 1692646696
transform 1 0 9568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1692646696
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1692646696
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1692646696
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_207
timestamp 1692646696
transform 1 0 20148 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_3
timestamp 1692646696
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_20
timestamp 1692646696
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1692646696
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_62
timestamp 1692646696
transform 1 0 6808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_74
timestamp 1692646696
transform 1 0 7912 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1692646696
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_98
timestamp 1692646696
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_115
timestamp 1692646696
transform 1 0 11684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_119
timestamp 1692646696
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_141
timestamp 1692646696
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_149
timestamp 1692646696
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_170
timestamp 1692646696
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_182
timestamp 1692646696
transform 1 0 17848 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_192
timestamp 1692646696
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1692646696
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_209
timestamp 1692646696
transform 1 0 20332 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_6
timestamp 1692646696
transform 1 0 1656 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_16
timestamp 1692646696
transform 1 0 2576 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_28
timestamp 1692646696
transform 1 0 3680 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_36
timestamp 1692646696
transform 1 0 4416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_48
timestamp 1692646696
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1692646696
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1692646696
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1692646696
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1692646696
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1692646696
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1692646696
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1692646696
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1692646696
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_137
timestamp 1692646696
transform 1 0 13708 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_144
timestamp 1692646696
transform 1 0 14352 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1692646696
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1692646696
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_173
timestamp 1692646696
transform 1 0 17020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_189
timestamp 1692646696
transform 1 0 18492 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_209
timestamp 1692646696
transform 1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1692646696
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1692646696
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_32
timestamp 1692646696
transform 1 0 4048 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1692646696
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1692646696
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1692646696
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_77
timestamp 1692646696
transform 1 0 8188 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 1692646696
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_88
timestamp 1692646696
transform 1 0 9200 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_97
timestamp 1692646696
transform 1 0 10028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_105
timestamp 1692646696
transform 1 0 10764 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_112
timestamp 1692646696
transform 1 0 11408 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_120
timestamp 1692646696
transform 1 0 12144 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_148
timestamp 1692646696
transform 1 0 14720 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_170
timestamp 1692646696
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1692646696
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1692646696
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_209
timestamp 1692646696
transform 1 0 20332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_3
timestamp 1692646696
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_15
timestamp 1692646696
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 1692646696
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_61
timestamp 1692646696
transform 1 0 6716 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_69
timestamp 1692646696
transform 1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_150
timestamp 1692646696
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_154
timestamp 1692646696
transform 1 0 15272 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_164
timestamp 1692646696
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1692646696
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_173
timestamp 1692646696
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_200
timestamp 1692646696
transform 1 0 19504 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_208
timestamp 1692646696
transform 1 0 20240 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_23
timestamp 1692646696
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp 1692646696
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_113
timestamp 1692646696
transform 1 0 11500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_125
timestamp 1692646696
transform 1 0 12604 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_133
timestamp 1692646696
transform 1 0 13340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_137
timestamp 1692646696
transform 1 0 13708 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_175
timestamp 1692646696
transform 1 0 17204 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1692646696
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_209
timestamp 1692646696
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_3
timestamp 1692646696
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_9
timestamp 1692646696
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_13
timestamp 1692646696
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_25
timestamp 1692646696
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_37
timestamp 1692646696
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_49
timestamp 1692646696
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1692646696
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_57
timestamp 1692646696
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_68
timestamp 1692646696
transform 1 0 7360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_80
timestamp 1692646696
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_89
timestamp 1692646696
transform 1 0 9292 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_95
timestamp 1692646696
transform 1 0 9844 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_100
timestamp 1692646696
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1692646696
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1692646696
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1692646696
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_137
timestamp 1692646696
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1692646696
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_186
timestamp 1692646696
transform 1 0 18216 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_208
timestamp 1692646696
transform 1 0 20240 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_23
timestamp 1692646696
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1692646696
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_49
timestamp 1692646696
transform 1 0 5612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_57
timestamp 1692646696
transform 1 0 6348 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_72
timestamp 1692646696
transform 1 0 7728 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_78
timestamp 1692646696
transform 1 0 8280 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1692646696
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1692646696
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_97
timestamp 1692646696
transform 1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_105
timestamp 1692646696
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_132
timestamp 1692646696
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp 1692646696
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_147
timestamp 1692646696
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_167
timestamp 1692646696
transform 1 0 16468 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_171
timestamp 1692646696
transform 1 0 16836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_183
timestamp 1692646696
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1692646696
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1692646696
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_209
timestamp 1692646696
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_3
timestamp 1692646696
transform 1 0 1380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_57
timestamp 1692646696
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_101
timestamp 1692646696
transform 1 0 10396 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_126
timestamp 1692646696
transform 1 0 12696 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_138
timestamp 1692646696
transform 1 0 13800 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_160
timestamp 1692646696
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_169
timestamp 1692646696
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_182
timestamp 1692646696
transform 1 0 17848 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_205
timestamp 1692646696
transform 1 0 19964 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1692646696
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1692646696
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1692646696
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_42
timestamp 1692646696
transform 1 0 4968 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_54
timestamp 1692646696
transform 1 0 6072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1692646696
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1692646696
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_85
timestamp 1692646696
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_108
timestamp 1692646696
transform 1 0 11040 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_135
timestamp 1692646696
transform 1 0 13524 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_163
timestamp 1692646696
transform 1 0 16100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_188
timestamp 1692646696
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_204
timestamp 1692646696
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_3
timestamp 1692646696
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_7
timestamp 1692646696
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_11
timestamp 1692646696
transform 1 0 2116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_23
timestamp 1692646696
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1692646696
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1692646696
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1692646696
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1692646696
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1692646696
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1692646696
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1692646696
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_93
timestamp 1692646696
transform 1 0 9660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_99
timestamp 1692646696
transform 1 0 10212 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_103
timestamp 1692646696
transform 1 0 10580 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1692646696
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1692646696
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_125
timestamp 1692646696
transform 1 0 12604 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_169
timestamp 1692646696
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_189
timestamp 1692646696
transform 1 0 18492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_210
timestamp 1692646696
transform 1 0 20424 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_7
timestamp 1692646696
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_38
timestamp 1692646696
transform 1 0 4600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_46
timestamp 1692646696
transform 1 0 5336 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_67
timestamp 1692646696
transform 1 0 7268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_79
timestamp 1692646696
transform 1 0 8372 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1692646696
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1692646696
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_97
timestamp 1692646696
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_123
timestamp 1692646696
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_135
timestamp 1692646696
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1692646696
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_141
timestamp 1692646696
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_162
timestamp 1692646696
transform 1 0 16008 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_174
timestamp 1692646696
transform 1 0 17112 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1692646696
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_209
timestamp 1692646696
transform 1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 1692646696
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_45
timestamp 1692646696
transform 1 0 5244 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_52
timestamp 1692646696
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1692646696
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_61
timestamp 1692646696
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1692646696
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1692646696
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_121
timestamp 1692646696
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_143
timestamp 1692646696
transform 1 0 14260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_155
timestamp 1692646696
transform 1 0 15364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_159
timestamp 1692646696
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1692646696
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_169
timestamp 1692646696
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_173
timestamp 1692646696
transform 1 0 17020 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_181
timestamp 1692646696
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_203
timestamp 1692646696
transform 1 0 19780 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_10
timestamp 1692646696
transform 1 0 2024 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_18
timestamp 1692646696
transform 1 0 2760 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_21
timestamp 1692646696
transform 1 0 3036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_25
timestamp 1692646696
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1692646696
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_72
timestamp 1692646696
transform 1 0 7728 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_80
timestamp 1692646696
transform 1 0 8464 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1692646696
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_103
timestamp 1692646696
transform 1 0 10580 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_115
timestamp 1692646696
transform 1 0 11684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_127
timestamp 1692646696
transform 1 0 12788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_135
timestamp 1692646696
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_158
timestamp 1692646696
transform 1 0 15640 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_176
timestamp 1692646696
transform 1 0 17296 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_187
timestamp 1692646696
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_191
timestamp 1692646696
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1692646696
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_204
timestamp 1692646696
transform 1 0 19872 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_210
timestamp 1692646696
transform 1 0 20424 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1692646696
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1692646696
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1692646696
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_42
timestamp 1692646696
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 1692646696
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_57
timestamp 1692646696
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_65
timestamp 1692646696
transform 1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_95
timestamp 1692646696
transform 1 0 9844 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_107
timestamp 1692646696
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1692646696
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_113
timestamp 1692646696
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_119
timestamp 1692646696
transform 1 0 12052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_162
timestamp 1692646696
transform 1 0 16008 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_203
timestamp 1692646696
transform 1 0 19780 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_3
timestamp 1692646696
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_21
timestamp 1692646696
transform 1 0 3036 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1692646696
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_29
timestamp 1692646696
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_44
timestamp 1692646696
transform 1 0 5152 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_52
timestamp 1692646696
transform 1 0 5888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_59
timestamp 1692646696
transform 1 0 6532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_63
timestamp 1692646696
transform 1 0 6900 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_71
timestamp 1692646696
transform 1 0 7636 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_75
timestamp 1692646696
transform 1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1692646696
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_88
timestamp 1692646696
transform 1 0 9200 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_100
timestamp 1692646696
transform 1 0 10304 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_108
timestamp 1692646696
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_129
timestamp 1692646696
transform 1 0 12972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1692646696
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_148
timestamp 1692646696
transform 1 0 14720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_152
timestamp 1692646696
transform 1 0 15088 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_177
timestamp 1692646696
transform 1 0 17388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_190
timestamp 1692646696
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_203
timestamp 1692646696
transform 1 0 19780 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1692646696
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_27
timestamp 1692646696
transform 1 0 3588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_74
timestamp 1692646696
transform 1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_99
timestamp 1692646696
transform 1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_103
timestamp 1692646696
transform 1 0 10580 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_130
timestamp 1692646696
transform 1 0 13064 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_152
timestamp 1692646696
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_164
timestamp 1692646696
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_169
timestamp 1692646696
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_177
timestamp 1692646696
transform 1 0 17388 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_187
timestamp 1692646696
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_191
timestamp 1692646696
transform 1 0 18676 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1692646696
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1692646696
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1692646696
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp 1692646696
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_35
timestamp 1692646696
transform 1 0 4324 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_47
timestamp 1692646696
transform 1 0 5428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_55
timestamp 1692646696
transform 1 0 6164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_59
timestamp 1692646696
transform 1 0 6532 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_68
timestamp 1692646696
transform 1 0 7360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_80
timestamp 1692646696
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1692646696
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_97
timestamp 1692646696
transform 1 0 10028 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_126
timestamp 1692646696
transform 1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_130
timestamp 1692646696
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1692646696
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_146
timestamp 1692646696
transform 1 0 14536 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_154
timestamp 1692646696
transform 1 0 15272 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_174
timestamp 1692646696
transform 1 0 17112 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1692646696
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_209
timestamp 1692646696
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1692646696
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1692646696
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_27
timestamp 1692646696
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_33
timestamp 1692646696
transform 1 0 4140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_42
timestamp 1692646696
transform 1 0 4968 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_50
timestamp 1692646696
transform 1 0 5704 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_81
timestamp 1692646696
transform 1 0 8556 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_85
timestamp 1692646696
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_97
timestamp 1692646696
transform 1 0 10028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_101
timestamp 1692646696
transform 1 0 10396 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_104
timestamp 1692646696
transform 1 0 10672 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_152
timestamp 1692646696
transform 1 0 15088 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_164
timestamp 1692646696
transform 1 0 16192 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_203
timestamp 1692646696
transform 1 0 19780 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1692646696
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1692646696
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1692646696
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1692646696
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_37
timestamp 1692646696
transform 1 0 4508 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_44
timestamp 1692646696
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_56
timestamp 1692646696
transform 1 0 6256 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_62
timestamp 1692646696
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_71
timestamp 1692646696
transform 1 0 7636 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_79
timestamp 1692646696
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_102
timestamp 1692646696
transform 1 0 10488 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_121
timestamp 1692646696
transform 1 0 12236 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_158
timestamp 1692646696
transform 1 0 15640 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_170
timestamp 1692646696
transform 1 0 16744 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1692646696
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1692646696
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_209
timestamp 1692646696
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1692646696
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_15
timestamp 1692646696
transform 1 0 2484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_23
timestamp 1692646696
transform 1 0 3220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_27
timestamp 1692646696
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_29
timestamp 1692646696
transform 1 0 3772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_41
timestamp 1692646696
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1692646696
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1692646696
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1692646696
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_81
timestamp 1692646696
transform 1 0 8556 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_85
timestamp 1692646696
transform 1 0 8924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_97
timestamp 1692646696
transform 1 0 10028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1692646696
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1692646696
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_123
timestamp 1692646696
transform 1 0 12420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_135
timestamp 1692646696
transform 1 0 13524 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_151
timestamp 1692646696
transform 1 0 14996 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_163
timestamp 1692646696
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1692646696
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1692646696
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_187
timestamp 1692646696
transform 1 0 18308 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_191
timestamp 1692646696
transform 1 0 18676 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_195
timestamp 1692646696
transform 1 0 19044 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_197
timestamp 1692646696
transform 1 0 19228 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_205
timestamp 1692646696
transform 1 0 19964 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 11224 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1692646696
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1692646696
transform -1 0 9108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 14076 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1692646696
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1692646696
transform -1 0 20516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1692646696
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1692646696
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1692646696
transform -1 0 19044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1692646696
transform 1 0 10396 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1692646696
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1692646696
transform 1 0 3312 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1692646696
transform -1 0 20516 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  output11
timestamp 1692646696
transform 1 0 20240 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1692646696
transform 1 0 20148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output13
timestamp 1692646696
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_36
timestamp 1692646696
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1692646696
transform -1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_37
timestamp 1692646696
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1692646696
transform -1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_38
timestamp 1692646696
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1692646696
transform -1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_39
timestamp 1692646696
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1692646696
transform -1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_40
timestamp 1692646696
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1692646696
transform -1 0 20792 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_41
timestamp 1692646696
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1692646696
transform -1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_42
timestamp 1692646696
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1692646696
transform -1 0 20792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_43
timestamp 1692646696
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1692646696
transform -1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_44
timestamp 1692646696
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1692646696
transform -1 0 20792 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_45
timestamp 1692646696
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1692646696
transform -1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_46
timestamp 1692646696
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1692646696
transform -1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_47
timestamp 1692646696
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1692646696
transform -1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_48
timestamp 1692646696
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1692646696
transform -1 0 20792 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_49
timestamp 1692646696
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1692646696
transform -1 0 20792 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_50
timestamp 1692646696
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1692646696
transform -1 0 20792 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_51
timestamp 1692646696
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1692646696
transform -1 0 20792 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_52
timestamp 1692646696
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1692646696
transform -1 0 20792 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_53
timestamp 1692646696
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1692646696
transform -1 0 20792 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_54
timestamp 1692646696
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1692646696
transform -1 0 20792 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_55
timestamp 1692646696
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1692646696
transform -1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_56
timestamp 1692646696
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1692646696
transform -1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_57
timestamp 1692646696
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1692646696
transform -1 0 20792 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_58
timestamp 1692646696
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1692646696
transform -1 0 20792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_59
timestamp 1692646696
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1692646696
transform -1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_60
timestamp 1692646696
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1692646696
transform -1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_61
timestamp 1692646696
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1692646696
transform -1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_62
timestamp 1692646696
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1692646696
transform -1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_63
timestamp 1692646696
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1692646696
transform -1 0 20792 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_64
timestamp 1692646696
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1692646696
transform -1 0 20792 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_65
timestamp 1692646696
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1692646696
transform -1 0 20792 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_66
timestamp 1692646696
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1692646696
transform -1 0 20792 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_67
timestamp 1692646696
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1692646696
transform -1 0 20792 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_68
timestamp 1692646696
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1692646696
transform -1 0 20792 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_69
timestamp 1692646696
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1692646696
transform -1 0 20792 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_70
timestamp 1692646696
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1692646696
transform -1 0 20792 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_71
timestamp 1692646696
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1692646696
transform -1 0 20792 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  PoR.ROSC_CLKBUF_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 2484 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  PoR.ROSC_CLKBUF_1
timestamp 1692646696
transform 1 0 1472 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYBUF_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 2392 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_0.clkdlybuf
timestamp 1692646696
transform -1 0 4968 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_0.clkinv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 5152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_1.clkdlybuf
timestamp 1692646696
transform 1 0 2484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_1.clkinv
timestamp 1692646696
transform -1 0 4324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_2.clkdlybuf
timestamp 1692646696
transform 1 0 1932 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_2.clkinv
timestamp 1692646696
transform 1 0 3220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_3.clkdlybuf
timestamp 1692646696
transform 1 0 1564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_3.clkinv
timestamp 1692646696
transform 1 0 2668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_4.clkdlybuf
timestamp 1692646696
transform -1 0 2300 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_4.clkinv
timestamp 1692646696
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_5.clkdlybuf
timestamp 1692646696
transform 1 0 1564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_5.clkinv
timestamp 1692646696
transform 1 0 1472 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  PoR.ROSC_DLYINV_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 2576 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1692646696
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1692646696
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1692646696
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1692646696
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1692646696
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1692646696
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1692646696
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1692646696
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1692646696
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_82
timestamp 1692646696
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_83
timestamp 1692646696
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1692646696
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1692646696
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_86
timestamp 1692646696
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_87
timestamp 1692646696
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_88
timestamp 1692646696
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_89
timestamp 1692646696
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_90
timestamp 1692646696
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_91
timestamp 1692646696
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_92
timestamp 1692646696
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_93
timestamp 1692646696
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_94
timestamp 1692646696
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_95
timestamp 1692646696
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_96
timestamp 1692646696
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_97
timestamp 1692646696
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_98
timestamp 1692646696
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_99
timestamp 1692646696
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_100
timestamp 1692646696
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_101
timestamp 1692646696
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp 1692646696
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_103
timestamp 1692646696
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_104
timestamp 1692646696
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_105
timestamp 1692646696
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_106
timestamp 1692646696
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_107
timestamp 1692646696
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_108
timestamp 1692646696
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp 1692646696
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_110
timestamp 1692646696
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_111
timestamp 1692646696
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp 1692646696
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp 1692646696
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp 1692646696
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp 1692646696
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp 1692646696
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_117
timestamp 1692646696
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_118
timestamp 1692646696
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_119
timestamp 1692646696
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_120
timestamp 1692646696
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_121
timestamp 1692646696
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_122
timestamp 1692646696
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_123
timestamp 1692646696
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_124
timestamp 1692646696
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_125
timestamp 1692646696
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_126
timestamp 1692646696
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_127
timestamp 1692646696
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_128
timestamp 1692646696
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_129
timestamp 1692646696
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_130
timestamp 1692646696
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_131
timestamp 1692646696
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_132
timestamp 1692646696
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_133
timestamp 1692646696
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_134
timestamp 1692646696
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_135
timestamp 1692646696
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_136
timestamp 1692646696
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_137
timestamp 1692646696
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_138
timestamp 1692646696
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_139
timestamp 1692646696
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_140
timestamp 1692646696
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_141
timestamp 1692646696
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_142
timestamp 1692646696
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_143
timestamp 1692646696
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_144
timestamp 1692646696
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_145
timestamp 1692646696
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_146
timestamp 1692646696
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_147
timestamp 1692646696
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_148
timestamp 1692646696
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_149
timestamp 1692646696
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_150
timestamp 1692646696
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_151
timestamp 1692646696
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_152
timestamp 1692646696
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_153
timestamp 1692646696
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_154
timestamp 1692646696
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_155
timestamp 1692646696
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_156
timestamp 1692646696
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_157
timestamp 1692646696
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_158
timestamp 1692646696
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_159
timestamp 1692646696
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_160
timestamp 1692646696
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_161
timestamp 1692646696
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_162
timestamp 1692646696
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_163
timestamp 1692646696
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_164
timestamp 1692646696
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_165
timestamp 1692646696
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_166
timestamp 1692646696
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_167
timestamp 1692646696
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_168
timestamp 1692646696
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_169
timestamp 1692646696
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_170
timestamp 1692646696
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_171
timestamp 1692646696
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_172
timestamp 1692646696
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_173
timestamp 1692646696
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_174
timestamp 1692646696
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_175
timestamp 1692646696
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_176
timestamp 1692646696
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_177
timestamp 1692646696
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_178
timestamp 1692646696
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_179
timestamp 1692646696
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_180
timestamp 1692646696
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_181
timestamp 1692646696
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_182
timestamp 1692646696
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_183
timestamp 1692646696
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_184
timestamp 1692646696
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_185
timestamp 1692646696
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_186
timestamp 1692646696
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_187
timestamp 1692646696
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_188
timestamp 1692646696
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_189
timestamp 1692646696
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_190
timestamp 1692646696
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1692646696
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1692646696
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1692646696
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_194
timestamp 1692646696
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_195
timestamp 1692646696
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_196
timestamp 1692646696
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_197
timestamp 1692646696
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_198
timestamp 1692646696
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_199
timestamp 1692646696
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_200
timestamp 1692646696
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_201
timestamp 1692646696
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_202
timestamp 1692646696
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_203
timestamp 1692646696
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_204
timestamp 1692646696
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
<< labels >>
flabel metal3 s 21118 15648 21918 15768 0 FreeSans 480 0 0 0 clk
port 0 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 clk_div[0]
port 1 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 clk_div[1]
port 2 nsew signal input
flabel metal2 s 13542 23262 13598 24062 0 FreeSans 224 90 0 0 one
port 3 nsew signal input
flabel metal2 s 8390 23262 8446 24062 0 FreeSans 224 90 0 0 por_fb_in
port 4 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 por_fb_out
port 5 nsew signal tristate
flabel metal3 s 21118 21088 21918 21208 0 FreeSans 480 0 0 0 por_n
port 6 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 rst_n
port 7 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 sel_mux0
port 8 nsew signal input
flabel metal3 s 21118 4768 21918 4888 0 FreeSans 480 0 0 0 sel_mux1
port 9 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 sel_mux2
port 10 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 sel_rosc[0]
port 11 nsew signal input
flabel metal2 s 18694 23262 18750 24062 0 FreeSans 224 90 0 0 sel_rosc[1]
port 12 nsew signal input
flabel metal4 s 4208 2128 4528 21808 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 10208 2128 10528 21808 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 16208 2128 16528 21808 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 7208 2128 7528 21808 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal4 s 13208 2128 13528 21808 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal4 s 19208 2128 19528 21808 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 xclk0
port 15 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 xclk1
port 16 nsew signal input
flabel metal2 s 3238 23262 3294 24062 0 FreeSans 224 90 0 0 xrst_n
port 17 nsew signal input
flabel metal3 s 21118 10208 21918 10328 0 FreeSans 480 0 0 0 zero
port 18 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 21918 24062
<< end >>
