/*
	Copyright 2020 Mohamed Shalan (mshalan@aucegypt.edu)
	
	Licensed under the Apache License, Version 2.0 (the "License"); 
	you may not use this file except in compliance with the License. 
	You may obtain a copy of the License at:
	http://www.apache.org/licenses/LICENSE-2.0
	Unless required by applicable law or agreed to in writing, software 
	distributed under the License is distributed on an "AS IS" BASIS, 
	WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
	See the License for the specific language governing permissions and 
	limitations under the License.
*/
/*
    All Digital Power-on-Reset (ADPoR) and Ring Oscillator (ROSC)
    (1) ADPoR
        - It asserts the rest (actibe low) for LENGTH clock cycles when the system is powered on.
        - Its clock is generated by a ring oscillator and is fixed @ 500KHz.
        - Assertion time is LENGTH x 2 micro-seconds
    (2) ROSC
        - A fixed clok output (8MHz)
        - A variable frequency clock output, 128/64/32/16 MHz (Selectable)
*/

`timescale          1ns/1ps
`default_nettype    none

module por_rosc #(parameter LENGTH=16) (
    input   wire        rst_n,          // System reset
    input   wire        fb_in,          // Oscillator feedback input
    input   wire        zero,           // Tie low 
    input   wire        one,            // Tie high 
    input   wire [1:0]  freq_sel,       // Select the frequency of clk_out; 0:128MHz, 1:64MHz, 2:32MHz, 3:16MHz
    output  wire        clk_8mhz,       // Fixed 8MHz clock
    output  wire        clk_128mhz,       // Fixed 128MHz clock
    output  wire        clk_out,        // Variable clock output; depends on freq_sel
    output  wire        por_n,          // Power on Reset output
    output  wire        fb_out          // Oscillator feedback output
);

`ifdef RTL_SIM
    reg         fake_clk = 0;
    assign      clk_128mhz = fake_clk;
    always #3.9 fake_clk = !fake_clk;
`else
    // 128MHz ROSC
    wire [8:1]  dly;
    //wire        clk_128mhz;

    (* keep *) sky130_fd_sc_hd__clkdlyinv5sd3_1    ROSC_DLYINV_0 ( .A(fb_in), .Y(dly[1]) );
    (* keep *) sky130_fd_sc_hd__clkdlyinv5sd3_1    ROSC_DLYINV_1 ( .A(dly[1]), .Y(dly[2]) );

    (* keep *) sky130_fd_sc_hd__clkdlyinv5sd3_1    ROSC_DLYINV_2 ( .A(dly[2]), .Y(dly[3]) );
    (* keep *) sky130_fd_sc_hd__clkdlyinv5sd3_1    ROSC_DLYINV_3 ( .A(dly[3]), .Y(dly[4]) );

    (* keep *) sky130_fd_sc_hd__clkdlyinv5sd3_1    ROSC_DLYINV_4 ( .A(dly[4]), .Y(dly[5]) );
    (* keep *) sky130_fd_sc_hd__clkdlyinv5sd3_1    ROSC_DLYINV_5 ( .A(dly[5]), .Y(dly[6]) );

    (* keep *) sky130_fd_sc_hd__clkdlybuf4s50_1    ROSC_DLYBUF_6 (.A(dly[6]), .X(dly[7]));
    
    (* keep *) sky130_fd_sc_hd__clkinv_8           ROSC_DLYINV_7 ( .A(dly[7]), .Y(dly[8]) );

    (* keep *) sky130_fd_sc_hd__clkbuf_8           ROSC_CLKBUF_0 ( .A(dly[8]), .X(fb_out) );
    (* keep *) sky130_fd_sc_hd__clkbuf_8           ROSC_CLKBUF_1 ( .A(fb_out), .X(clk_128mhz) );

`endif
    // Clock Divider
    (* keep *) reg [8:1]   clk_div = 0;    // The initialization is needed only for simulation
    wire        clk_64mhz  = clk_div[1];
    wire        clk_32mhz  = clk_div[2];
    wire        clk_16mhz  = clk_div[3];
    wire        clk_500khz = clk_div[8];
    
    assign      clk_8mhz   = clk_div[4];

    (* keep *)
    always @(posedge clk_128mhz)
        clk_div <= clk_div + 1'b1;
    
    // Frequency 4x1 MUX
    clkmux_4x1 CLKMUX (
        .rst_n(rst_n),
        .clk1(clk_128mhz), 
        .clk2(clk_64mhz), 
        .clk3(clk_32mhz), 
        .clk4(clk_16mhz),
        .sel(freq_sel),
        .clko(clk_out)
    );
    
    // All digital PoR
`ifdef RTL_SIM
    (* keep *) reg [LENGTH-1:0] shift_reg0 = 16'hDEAD;
    (* keep *) reg [LENGTH-1:0] shift_reg1 = 16'hBEEF;
    (* keep *) reg [LENGTH-1:0] shift_reg2 = 16'hDEAF;
    (* keep *) reg [LENGTH-1:0] shift_reg3 = 16'hBEAD;
`else
    (* keep *) reg [LENGTH-1:0] shift_reg0;
    (* keep *) reg [LENGTH-1:0] shift_reg1;
    (* keep *) reg [LENGTH-1:0] shift_reg2;
    (* keep *) reg [LENGTH-1:0] shift_reg3;
`endif

    (* keep *)
    wire cmp0, cmp1, cmp2, cmp3;

    (* keep *)
    always @(posedge clk_500khz) begin
        (* keep *) shift_reg0 <= {one, shift_reg0[LENGTH-1:1]};
        (* keep *) shift_reg1 <= {zero, shift_reg1[LENGTH-1:1]};
        (* keep *) shift_reg2 <= {one, shift_reg2[LENGTH-1:1]};
        (* keep *) shift_reg3 <= {zero, shift_reg3[LENGTH-1:1]};
    end

    assign cmp0 = (shift_reg0 == {LENGTH{one}});
    assign cmp1 = (shift_reg1 == {LENGTH{zero}});
    assign cmp2 = (shift_reg2 == {LENGTH{one}});
    assign cmp3 = (shift_reg3 == {LENGTH{zero}});

    assign por_n = cmp0 & cmp1 & cmp2 & cmp3;    


endmodule

`ifndef RTL_SIM
module sky130_fd_sc_hd__clkdlyinv5sd3_1 (output Y, input  A);
    // Local signals
    wire clkinv_out;
    // Mapping
    sky130_fd_sc_hd__clkinv_2 clkinv (
        .A(A), 
        .Y(clkinv_out)
    );
    sky130_fd_sc_hd__clkdlybuf4s50_1 clkdlybuf (
        .A(clkinv_out), 
        .X(Y)
    );
endmodule
`endif