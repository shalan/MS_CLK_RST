magic
tech sky130A
magscale 1 2
timestamp 1693235701
<< viali >>
rect 1409 17629 1443 17663
rect 2881 17629 2915 17663
rect 16129 17629 16163 17663
rect 16405 17629 16439 17663
rect 1593 17493 1627 17527
rect 2697 17493 2731 17527
rect 15945 17493 15979 17527
rect 16221 17493 16255 17527
rect 2421 17153 2455 17187
rect 6193 17153 6227 17187
rect 10425 17153 10459 17187
rect 10701 17153 10735 17187
rect 11161 17153 11195 17187
rect 2697 17085 2731 17119
rect 11529 17085 11563 17119
rect 11805 17085 11839 17119
rect 13369 17085 13403 17119
rect 13737 17017 13771 17051
rect 4169 16949 4203 16983
rect 5549 16949 5583 16983
rect 11253 16949 11287 16983
rect 13277 16949 13311 16983
rect 13829 16949 13863 16983
rect 2789 16745 2823 16779
rect 11345 16745 11379 16779
rect 2605 16677 2639 16711
rect 4077 16609 4111 16643
rect 11713 16609 11747 16643
rect 11989 16609 12023 16643
rect 2881 16541 2915 16575
rect 2973 16541 3007 16575
rect 3801 16541 3835 16575
rect 5641 16541 5675 16575
rect 11345 16541 11379 16575
rect 11529 16541 11563 16575
rect 13737 16541 13771 16575
rect 14197 16541 14231 16575
rect 2329 16473 2363 16507
rect 5549 16405 5583 16439
rect 5825 16405 5859 16439
rect 13461 16405 13495 16439
rect 13553 16405 13587 16439
rect 14289 16405 14323 16439
rect 12909 16133 12943 16167
rect 13553 16133 13587 16167
rect 1409 16065 1443 16099
rect 1869 16065 1903 16099
rect 1961 16065 1995 16099
rect 2053 16065 2087 16099
rect 2237 16065 2271 16099
rect 2421 16065 2455 16099
rect 2697 16065 2731 16099
rect 2881 16065 2915 16099
rect 5917 16065 5951 16099
rect 12725 16065 12759 16099
rect 12817 16065 12851 16099
rect 13093 16065 13127 16099
rect 13277 15997 13311 16031
rect 1593 15929 1627 15963
rect 2513 15929 2547 15963
rect 1685 15861 1719 15895
rect 2697 15861 2731 15895
rect 5273 15861 5307 15895
rect 12541 15861 12575 15895
rect 15025 15861 15059 15895
rect 5812 15657 5846 15691
rect 8585 15657 8619 15691
rect 9321 15589 9355 15623
rect 14381 15589 14415 15623
rect 1777 15521 1811 15555
rect 2053 15521 2087 15555
rect 5549 15521 5583 15555
rect 9413 15521 9447 15555
rect 15853 15521 15887 15555
rect 16129 15521 16163 15555
rect 5457 15453 5491 15487
rect 8585 15453 8619 15487
rect 8769 15453 8803 15487
rect 9689 15453 9723 15487
rect 9873 15453 9907 15487
rect 4721 15385 4755 15419
rect 8953 15385 8987 15419
rect 3525 15317 3559 15351
rect 4813 15317 4847 15351
rect 7297 15317 7331 15351
rect 8493 15317 8527 15351
rect 9505 15317 9539 15351
rect 9965 15317 9999 15351
rect 11437 15317 11471 15351
rect 5365 15113 5399 15147
rect 8677 15113 8711 15147
rect 9597 15113 9631 15147
rect 13261 15113 13295 15147
rect 2237 15045 2271 15079
rect 3065 15045 3099 15079
rect 7205 15045 7239 15079
rect 9137 15045 9171 15079
rect 13461 15045 13495 15079
rect 13645 15045 13679 15079
rect 13829 15045 13863 15079
rect 1961 14977 1995 15011
rect 2145 14977 2179 15011
rect 2329 14977 2363 15011
rect 2789 14977 2823 15011
rect 4813 14977 4847 15011
rect 5365 14977 5399 15011
rect 6193 14977 6227 15011
rect 6653 14977 6687 15011
rect 8861 14977 8895 15011
rect 9045 14977 9079 15011
rect 9234 14977 9268 15011
rect 11529 14977 11563 15011
rect 11785 14977 11819 15011
rect 13553 14977 13587 15011
rect 15393 14977 15427 15011
rect 4537 14909 4571 14943
rect 6745 14909 6779 14943
rect 6929 14909 6963 14943
rect 11069 14909 11103 14943
rect 11345 14909 11379 14943
rect 15301 14909 15335 14943
rect 2513 14773 2547 14807
rect 4813 14773 4847 14807
rect 9413 14773 9447 14807
rect 12909 14773 12943 14807
rect 13093 14773 13127 14807
rect 13277 14773 13311 14807
rect 13829 14773 13863 14807
rect 15669 14773 15703 14807
rect 7021 14569 7055 14603
rect 10701 14569 10735 14603
rect 12265 14569 12299 14603
rect 13829 14569 13863 14603
rect 16681 14501 16715 14535
rect 7113 14433 7147 14467
rect 9229 14433 9263 14467
rect 11161 14433 11195 14467
rect 11437 14433 11471 14467
rect 4629 14365 4663 14399
rect 8953 14365 8987 14399
rect 11069 14365 11103 14399
rect 12449 14365 12483 14399
rect 15301 14365 15335 14399
rect 15568 14365 15602 14399
rect 7380 14297 7414 14331
rect 12716 14297 12750 14331
rect 3985 14229 4019 14263
rect 8493 14229 8527 14263
rect 15117 14229 15151 14263
rect 7849 14025 7883 14059
rect 13093 14025 13127 14059
rect 15393 14025 15427 14059
rect 15761 13957 15795 13991
rect 4077 13889 4111 13923
rect 4169 13889 4203 13923
rect 7941 13889 7975 13923
rect 10057 13889 10091 13923
rect 13001 13889 13035 13923
rect 13185 13889 13219 13923
rect 14280 13889 14314 13923
rect 15945 13889 15979 13923
rect 4445 13821 4479 13855
rect 10149 13821 10183 13855
rect 14013 13821 14047 13855
rect 3433 13685 3467 13719
rect 13921 13685 13955 13719
rect 15577 13685 15611 13719
rect 14657 13481 14691 13515
rect 15577 13481 15611 13515
rect 9137 13345 9171 13379
rect 12081 13345 12115 13379
rect 15393 13345 15427 13379
rect 3433 13277 3467 13311
rect 6285 13277 6319 13311
rect 13829 13277 13863 13311
rect 14841 13277 14875 13311
rect 15025 13277 15059 13311
rect 15209 13277 15243 13311
rect 15485 13277 15519 13311
rect 15669 13277 15703 13311
rect 6561 13209 6595 13243
rect 9413 13209 9447 13243
rect 13553 13209 13587 13243
rect 3433 13141 3467 13175
rect 8033 13141 8067 13175
rect 10885 13141 10919 13175
rect 7205 12937 7239 12971
rect 9321 12937 9355 12971
rect 10701 12937 10735 12971
rect 10977 12937 11011 12971
rect 13277 12937 13311 12971
rect 2697 12869 2731 12903
rect 7665 12869 7699 12903
rect 9965 12869 9999 12903
rect 11805 12869 11839 12903
rect 15117 12869 15151 12903
rect 15317 12869 15351 12903
rect 2881 12801 2915 12835
rect 3157 12801 3191 12835
rect 4997 12801 5031 12835
rect 5641 12801 5675 12835
rect 7113 12801 7147 12835
rect 7389 12801 7423 12835
rect 9229 12801 9263 12835
rect 9413 12801 9447 12835
rect 9729 12801 9763 12835
rect 9873 12801 9907 12835
rect 10149 12801 10183 12835
rect 10793 12801 10827 12835
rect 11529 12801 11563 12835
rect 16313 12801 16347 12835
rect 5733 12733 5767 12767
rect 6929 12733 6963 12767
rect 10241 12733 10275 12767
rect 5273 12665 5307 12699
rect 6653 12665 6687 12699
rect 9597 12665 9631 12699
rect 10609 12665 10643 12699
rect 3065 12597 3099 12631
rect 4813 12597 4847 12631
rect 6469 12597 6503 12631
rect 9137 12597 9171 12631
rect 14289 12597 14323 12631
rect 15301 12597 15335 12631
rect 15485 12597 15519 12631
rect 16497 12597 16531 12631
rect 6653 12393 6687 12427
rect 12265 12393 12299 12427
rect 12449 12393 12483 12427
rect 14381 12393 14415 12427
rect 6101 12325 6135 12359
rect 1869 12257 1903 12291
rect 10517 12257 10551 12291
rect 10793 12257 10827 12291
rect 4721 12189 4755 12223
rect 4988 12189 5022 12223
rect 6837 12189 6871 12223
rect 12541 12189 12575 12223
rect 13369 12189 13403 12223
rect 13553 12189 13587 12223
rect 14105 12189 14139 12223
rect 14197 12189 14231 12223
rect 15945 12189 15979 12223
rect 16037 12189 16071 12223
rect 16221 12189 16255 12223
rect 2145 12121 2179 12155
rect 13737 12121 13771 12155
rect 14381 12121 14415 12155
rect 15700 12121 15734 12155
rect 16129 12121 16163 12155
rect 3617 12053 3651 12087
rect 14565 12053 14599 12087
rect 5281 11849 5315 11883
rect 14381 11849 14415 11883
rect 3157 11781 3191 11815
rect 7573 11781 7607 11815
rect 9689 11781 9723 11815
rect 14841 11781 14875 11815
rect 2881 11713 2915 11747
rect 4721 11713 4755 11747
rect 4905 11713 4939 11747
rect 4997 11713 5031 11747
rect 5094 11713 5128 11747
rect 7021 11713 7055 11747
rect 7205 11713 7239 11747
rect 7389 11713 7423 11747
rect 7665 11713 7699 11747
rect 7757 11713 7791 11747
rect 10885 11713 10919 11747
rect 12725 11713 12759 11747
rect 12909 11713 12943 11747
rect 13268 11713 13302 11747
rect 15025 11713 15059 11747
rect 15292 11713 15326 11747
rect 13001 11645 13035 11679
rect 4629 11509 4663 11543
rect 7021 11509 7055 11543
rect 7941 11509 7975 11543
rect 9413 11509 9447 11543
rect 10977 11509 11011 11543
rect 12541 11509 12575 11543
rect 12909 11509 12943 11543
rect 16405 11509 16439 11543
rect 2605 11305 2639 11339
rect 13553 11305 13587 11339
rect 15485 11305 15519 11339
rect 4629 11237 4663 11271
rect 6193 11169 6227 11203
rect 6377 11169 6411 11203
rect 7205 11169 7239 11203
rect 9873 11169 9907 11203
rect 11621 11169 11655 11203
rect 11989 11169 12023 11203
rect 15025 11169 15059 11203
rect 2421 11101 2455 11135
rect 2605 11101 2639 11135
rect 4077 11101 4111 11135
rect 4497 11101 4531 11135
rect 6009 11101 6043 11135
rect 6285 11101 6319 11135
rect 6469 11101 6503 11135
rect 6929 11101 6963 11135
rect 11713 11101 11747 11135
rect 13553 11101 13587 11135
rect 13737 11101 13771 11135
rect 15117 11101 15151 11135
rect 4261 11033 4295 11067
rect 4353 11033 4387 11067
rect 10149 11033 10183 11067
rect 5825 10965 5859 10999
rect 8677 10965 8711 10999
rect 13461 10965 13495 10999
rect 6377 10761 6411 10795
rect 9873 10761 9907 10795
rect 10517 10761 10551 10795
rect 3065 10693 3099 10727
rect 6745 10693 6779 10727
rect 8401 10693 8435 10727
rect 15025 10693 15059 10727
rect 2789 10625 2823 10659
rect 2973 10625 3007 10659
rect 3209 10625 3243 10659
rect 4813 10625 4847 10659
rect 5080 10625 5114 10659
rect 6561 10625 6595 10659
rect 7757 10625 7791 10659
rect 10701 10625 10735 10659
rect 12909 10625 12943 10659
rect 14289 10625 14323 10659
rect 14841 10625 14875 10659
rect 15117 10625 15151 10659
rect 15214 10625 15248 10659
rect 1409 10557 1443 10591
rect 7849 10557 7883 10591
rect 8125 10557 8159 10591
rect 10793 10557 10827 10591
rect 11253 10557 11287 10591
rect 13185 10557 13219 10591
rect 14013 10557 14047 10591
rect 6193 10489 6227 10523
rect 10977 10489 11011 10523
rect 15393 10489 15427 10523
rect 3341 10421 3375 10455
rect 13369 10421 13403 10455
rect 14197 10421 14231 10455
rect 3525 10217 3559 10251
rect 5549 10217 5583 10251
rect 14289 10217 14323 10251
rect 4629 10149 4663 10183
rect 11345 10149 11379 10183
rect 1593 10081 1627 10115
rect 11989 10081 12023 10115
rect 16497 10081 16531 10115
rect 3617 10013 3651 10047
rect 4077 10013 4111 10047
rect 4497 10013 4531 10047
rect 5733 10013 5767 10047
rect 6285 10013 6319 10047
rect 6377 10013 6411 10047
rect 10793 10013 10827 10047
rect 11069 10013 11103 10047
rect 11166 10013 11200 10047
rect 11529 10013 11563 10047
rect 11713 10013 11747 10047
rect 16773 10013 16807 10047
rect 1869 9945 1903 9979
rect 4261 9945 4295 9979
rect 4353 9945 4387 9979
rect 6193 9945 6227 9979
rect 6622 9945 6656 9979
rect 10977 9945 11011 9979
rect 12265 9945 12299 9979
rect 14197 9945 14231 9979
rect 3341 9877 3375 9911
rect 7757 9877 7791 9911
rect 11621 9877 11655 9911
rect 13737 9877 13771 9911
rect 15025 9877 15059 9911
rect 1961 9673 1995 9707
rect 4537 9673 4571 9707
rect 11253 9673 11287 9707
rect 11897 9673 11931 9707
rect 14933 9673 14967 9707
rect 13001 9605 13035 9639
rect 15393 9605 15427 9639
rect 1869 9537 1903 9571
rect 2053 9537 2087 9571
rect 2789 9537 2823 9571
rect 4813 9537 4847 9571
rect 11713 9537 11747 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 13185 9537 13219 9571
rect 15025 9537 15059 9571
rect 15209 9537 15243 9571
rect 15477 9537 15511 9571
rect 3065 9469 3099 9503
rect 7665 9469 7699 9503
rect 7941 9469 7975 9503
rect 9505 9469 9539 9503
rect 9781 9469 9815 9503
rect 13461 9469 13495 9503
rect 9413 9401 9447 9435
rect 4997 9333 5031 9367
rect 15025 9333 15059 9367
rect 2145 9129 2179 9163
rect 9505 9129 9539 9163
rect 11437 9129 11471 9163
rect 13921 9129 13955 9163
rect 16129 9129 16163 9163
rect 7113 9061 7147 9095
rect 4537 8993 4571 9027
rect 4721 8993 4755 9027
rect 13369 8993 13403 9027
rect 14657 8993 14691 9027
rect 2053 8925 2087 8959
rect 4629 8925 4663 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 6837 8925 6871 8959
rect 6981 8925 7015 8959
rect 7665 8925 7699 8959
rect 9413 8925 9447 8959
rect 14289 8925 14323 8959
rect 14381 8925 14415 8959
rect 4997 8857 5031 8891
rect 14197 8857 14231 8891
rect 6469 8789 6503 8823
rect 7757 8789 7791 8823
rect 5181 8585 5215 8619
rect 6377 8517 6411 8551
rect 8125 8517 8159 8551
rect 11345 8517 11379 8551
rect 13001 8517 13035 8551
rect 3433 8449 3467 8483
rect 5825 8449 5859 8483
rect 6009 8449 6043 8483
rect 7113 8449 7147 8483
rect 7849 8449 7883 8483
rect 11161 8449 11195 8483
rect 11529 8449 11563 8483
rect 11785 8449 11819 8483
rect 13277 8449 13311 8483
rect 13461 8449 13495 8483
rect 13553 8449 13587 8483
rect 13737 8449 13771 8483
rect 13921 8449 13955 8483
rect 16497 8449 16531 8483
rect 3709 8381 3743 8415
rect 5917 8381 5951 8415
rect 6837 8381 6871 8415
rect 9597 8381 9631 8415
rect 16221 8381 16255 8415
rect 6653 8313 6687 8347
rect 10977 8313 11011 8347
rect 12909 8313 12943 8347
rect 13369 8313 13403 8347
rect 6929 8245 6963 8279
rect 14565 8245 14599 8279
rect 14749 8245 14783 8279
rect 8401 8041 8435 8075
rect 10885 8041 10919 8075
rect 11621 8041 11655 8075
rect 13277 8041 13311 8075
rect 6653 7905 6687 7939
rect 6929 7905 6963 7939
rect 14105 7905 14139 7939
rect 3433 7837 3467 7871
rect 9413 7837 9447 7871
rect 9505 7837 9539 7871
rect 11437 7837 11471 7871
rect 13461 7837 13495 7871
rect 13553 7837 13587 7871
rect 13737 7837 13771 7871
rect 13829 7837 13863 7871
rect 9772 7769 9806 7803
rect 13185 7769 13219 7803
rect 14381 7769 14415 7803
rect 2789 7701 2823 7735
rect 15853 7701 15887 7735
rect 9781 7497 9815 7531
rect 11805 7497 11839 7531
rect 13737 7497 13771 7531
rect 14749 7497 14783 7531
rect 4445 7429 4479 7463
rect 9321 7429 9355 7463
rect 14197 7429 14231 7463
rect 16221 7429 16255 7463
rect 2973 7361 3007 7395
rect 9505 7361 9539 7395
rect 9689 7361 9723 7395
rect 9965 7361 9999 7395
rect 11989 7361 12023 7395
rect 16497 7361 16531 7395
rect 4169 7293 4203 7327
rect 12265 7293 12299 7327
rect 3617 7157 3651 7191
rect 4077 7157 4111 7191
rect 5917 7157 5951 7191
rect 13921 7157 13955 7191
rect 5996 6953 6030 6987
rect 9321 6953 9355 6987
rect 13369 6953 13403 6987
rect 16589 6953 16623 6987
rect 9873 6885 9907 6919
rect 12909 6885 12943 6919
rect 7573 6817 7607 6851
rect 8033 6817 8067 6851
rect 10149 6817 10183 6851
rect 12173 6817 12207 6851
rect 12265 6817 12299 6851
rect 12357 6817 12391 6851
rect 12450 6817 12484 6851
rect 5733 6749 5767 6783
rect 7941 6749 7975 6783
rect 8953 6749 8987 6783
rect 9597 6749 9631 6783
rect 9689 6749 9723 6783
rect 10057 6749 10091 6783
rect 12633 6749 12667 6783
rect 12909 6749 12943 6783
rect 16773 6749 16807 6783
rect 10425 6681 10459 6715
rect 13277 6681 13311 6715
rect 5641 6613 5675 6647
rect 7481 6613 7515 6647
rect 9321 6613 9355 6647
rect 9505 6613 9539 6647
rect 11897 6613 11931 6647
rect 11989 6613 12023 6647
rect 12725 6613 12759 6647
rect 8769 6409 8803 6443
rect 10057 6409 10091 6443
rect 10609 6409 10643 6443
rect 12081 6409 12115 6443
rect 13829 6409 13863 6443
rect 14197 6341 14231 6375
rect 3617 6273 3651 6307
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 4988 6273 5022 6307
rect 7297 6273 7331 6307
rect 7389 6273 7423 6307
rect 7656 6273 7690 6307
rect 10793 6273 10827 6307
rect 11989 6273 12023 6307
rect 12173 6273 12207 6307
rect 13645 6273 13679 6307
rect 2697 6205 2731 6239
rect 13921 6205 13955 6239
rect 13553 6137 13587 6171
rect 6101 6069 6135 6103
rect 15669 6069 15703 6103
rect 4905 5865 4939 5899
rect 10885 5865 10919 5899
rect 11161 5865 11195 5899
rect 14105 5865 14139 5899
rect 4629 5729 4663 5763
rect 10517 5729 10551 5763
rect 11805 5729 11839 5763
rect 14749 5729 14783 5763
rect 2697 5661 2731 5695
rect 4537 5661 4571 5695
rect 9781 5661 9815 5695
rect 9965 5661 9999 5695
rect 10057 5661 10091 5695
rect 11529 5661 11563 5695
rect 12725 5661 12759 5695
rect 12909 5661 12943 5695
rect 14473 5661 14507 5695
rect 14933 5661 14967 5695
rect 3433 5593 3467 5627
rect 10425 5593 10459 5627
rect 10885 5593 10919 5627
rect 13921 5593 13955 5627
rect 15209 5593 15243 5627
rect 5181 5525 5215 5559
rect 7757 5525 7791 5559
rect 11069 5525 11103 5559
rect 11621 5525 11655 5559
rect 12817 5525 12851 5559
rect 14565 5525 14599 5559
rect 16681 5525 16715 5559
rect 1593 5321 1627 5355
rect 4905 5321 4939 5355
rect 11805 5321 11839 5355
rect 14289 5321 14323 5355
rect 5273 5253 5307 5287
rect 5549 5253 5583 5287
rect 5749 5253 5783 5287
rect 8125 5253 8159 5287
rect 11253 5253 11287 5287
rect 12081 5253 12115 5287
rect 12633 5253 12667 5287
rect 14565 5253 14599 5287
rect 1409 5185 1443 5219
rect 3792 5185 3826 5219
rect 5181 5185 5215 5219
rect 5457 5185 5491 5219
rect 7021 5185 7055 5219
rect 7849 5185 7883 5219
rect 11161 5185 11195 5219
rect 11345 5185 11379 5219
rect 11713 5185 11747 5219
rect 11897 5185 11931 5219
rect 12449 5185 12483 5219
rect 13645 5185 13679 5219
rect 13803 5185 13837 5219
rect 13921 5185 13955 5219
rect 14013 5185 14047 5219
rect 14105 5185 14139 5219
rect 14749 5185 14783 5219
rect 14841 5185 14875 5219
rect 15025 5185 15059 5219
rect 3525 5117 3559 5151
rect 7297 5117 7331 5151
rect 7757 5117 7791 5151
rect 9597 5117 9631 5151
rect 7481 5049 7515 5083
rect 11529 5049 11563 5083
rect 14381 5049 14415 5083
rect 5457 4981 5491 5015
rect 5733 4981 5767 5015
rect 5917 4981 5951 5015
rect 7205 4981 7239 5015
rect 12265 4981 12299 5015
rect 14933 4981 14967 5015
rect 4169 4777 4203 4811
rect 9229 4777 9263 4811
rect 12725 4777 12759 4811
rect 13369 4777 13403 4811
rect 13553 4777 13587 4811
rect 14289 4777 14323 4811
rect 11161 4709 11195 4743
rect 11897 4709 11931 4743
rect 4997 4641 5031 4675
rect 9321 4641 9355 4675
rect 9597 4641 9631 4675
rect 11805 4641 11839 4675
rect 12081 4641 12115 4675
rect 12633 4641 12667 4675
rect 13277 4641 13311 4675
rect 4261 4573 4295 4607
rect 5089 4573 5123 4607
rect 5273 4573 5307 4607
rect 5365 4573 5399 4607
rect 7113 4573 7147 4607
rect 11345 4573 11379 4607
rect 11437 4573 11471 4607
rect 12173 4573 12207 4607
rect 12265 4573 12299 4607
rect 12357 4573 12391 4607
rect 12541 4573 12575 4607
rect 12817 4573 12851 4607
rect 13369 4573 13403 4607
rect 5181 4505 5215 4539
rect 5610 4505 5644 4539
rect 7358 4505 7392 4539
rect 11713 4505 11747 4539
rect 13093 4505 13127 4539
rect 14473 4505 14507 4539
rect 6745 4437 6779 4471
rect 8493 4437 8527 4471
rect 11069 4437 11103 4471
rect 13001 4437 13035 4471
rect 14105 4437 14139 4471
rect 14273 4437 14307 4471
rect 14749 4437 14783 4471
rect 5825 4233 5859 4267
rect 6009 4233 6043 4267
rect 7021 4233 7055 4267
rect 7481 4233 7515 4267
rect 8309 4233 8343 4267
rect 8401 4233 8435 4267
rect 11069 4233 11103 4267
rect 3249 4165 3283 4199
rect 4077 4165 4111 4199
rect 5641 4165 5675 4199
rect 5917 4165 5951 4199
rect 8125 4165 8159 4199
rect 13737 4165 13771 4199
rect 13921 4165 13955 4199
rect 14105 4165 14139 4199
rect 6377 4097 6411 4131
rect 6561 4097 6595 4131
rect 7941 4097 7975 4131
rect 8493 4097 8527 4131
rect 10885 4097 10919 4131
rect 11069 4097 11103 4131
rect 12633 4097 12667 4131
rect 12817 4097 12851 4131
rect 13277 4097 13311 4131
rect 13461 4097 13495 4131
rect 14381 4097 14415 4131
rect 14473 4097 14507 4131
rect 14749 4097 14783 4131
rect 7665 4029 7699 4063
rect 7757 4029 7791 4063
rect 7849 4029 7883 4063
rect 8677 4029 8711 4063
rect 13369 4029 13403 4063
rect 14013 4029 14047 4063
rect 15025 4029 15059 4063
rect 6193 3961 6227 3995
rect 13553 3961 13587 3995
rect 14657 3961 14691 3995
rect 6377 3893 6411 3927
rect 12817 3893 12851 3927
rect 16497 3893 16531 3927
rect 4813 3689 4847 3723
rect 6285 3689 6319 3723
rect 13185 3689 13219 3723
rect 4905 3553 4939 3587
rect 6377 3485 6411 3519
rect 6561 3485 6595 3519
rect 7665 3485 7699 3519
rect 7849 3485 7883 3519
rect 8033 3485 8067 3519
rect 8309 3485 8343 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 8769 3485 8803 3519
rect 11069 3485 11103 3519
rect 11161 3485 11195 3519
rect 11437 3485 11471 3519
rect 11529 3485 11563 3519
rect 11713 3485 11747 3519
rect 12449 3485 12483 3519
rect 12909 3485 12943 3519
rect 13461 3485 13495 3519
rect 13645 3485 13679 3519
rect 14105 3485 14139 3519
rect 14381 3485 14415 3519
rect 14473 3485 14507 3519
rect 5172 3417 5206 3451
rect 6469 3417 6503 3451
rect 8677 3417 8711 3451
rect 11253 3417 11287 3451
rect 11621 3417 11655 3451
rect 12541 3417 12575 3451
rect 12633 3417 12667 3451
rect 12751 3417 12785 3451
rect 13369 3417 13403 3451
rect 14289 3417 14323 3451
rect 8125 3349 8159 3383
rect 10885 3349 10919 3383
rect 12265 3349 12299 3383
rect 13001 3349 13035 3383
rect 13169 3349 13203 3383
rect 13829 3349 13863 3383
rect 14657 3349 14691 3383
rect 8033 3145 8067 3179
rect 13645 3145 13679 3179
rect 6193 3077 6227 3111
rect 9873 3077 9907 3111
rect 11805 3077 11839 3111
rect 13829 3077 13863 3111
rect 15577 3077 15611 3111
rect 6653 3009 6687 3043
rect 6920 3009 6954 3043
rect 9238 3009 9272 3043
rect 9505 3009 9539 3043
rect 9597 3009 9631 3043
rect 11529 3009 11563 3043
rect 13737 3009 13771 3043
rect 13921 3009 13955 3043
rect 15853 3009 15887 3043
rect 13277 2941 13311 2975
rect 14105 2941 14139 2975
rect 11345 2873 11379 2907
rect 8125 2805 8159 2839
rect 7205 2601 7239 2635
rect 7849 2601 7883 2635
rect 9505 2601 9539 2635
rect 9965 2601 9999 2635
rect 11713 2601 11747 2635
rect 16313 2601 16347 2635
rect 8493 2533 8527 2567
rect 8217 2465 8251 2499
rect 4813 2397 4847 2431
rect 7389 2397 7423 2431
rect 8125 2397 8159 2431
rect 9781 2397 9815 2431
rect 16497 2397 16531 2431
rect 4629 2329 4663 2363
<< metal1 >>
rect 1104 17978 17112 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 10214 17978
rect 10266 17926 10278 17978
rect 10330 17926 10342 17978
rect 10394 17926 10406 17978
rect 10458 17926 10470 17978
rect 10522 17926 16214 17978
rect 16266 17926 16278 17978
rect 16330 17926 16342 17978
rect 16394 17926 16406 17978
rect 16458 17926 16470 17978
rect 16522 17926 17112 17978
rect 1104 17904 17112 17926
rect 658 17688 664 17740
rect 716 17728 722 17740
rect 17034 17728 17040 17740
rect 716 17700 1440 17728
rect 716 17688 722 17700
rect 1412 17669 1440 17700
rect 16132 17700 17040 17728
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 2866 17620 2872 17672
rect 2924 17620 2930 17672
rect 16132 17669 16160 17700
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 16117 17663 16175 17669
rect 16117 17629 16129 17663
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 16206 17620 16212 17672
rect 16264 17660 16270 17672
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 16264 17632 16405 17660
rect 16264 17620 16270 17632
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 1578 17484 1584 17536
rect 1636 17484 1642 17536
rect 2682 17484 2688 17536
rect 2740 17484 2746 17536
rect 15930 17484 15936 17536
rect 15988 17484 15994 17536
rect 16206 17484 16212 17536
rect 16264 17484 16270 17536
rect 1104 17434 17112 17456
rect 1104 17382 7214 17434
rect 7266 17382 7278 17434
rect 7330 17382 7342 17434
rect 7394 17382 7406 17434
rect 7458 17382 7470 17434
rect 7522 17382 13214 17434
rect 13266 17382 13278 17434
rect 13330 17382 13342 17434
rect 13394 17382 13406 17434
rect 13458 17382 13470 17434
rect 13522 17382 17112 17434
rect 1104 17360 17112 17382
rect 2590 17280 2596 17332
rect 2648 17320 2654 17332
rect 15930 17320 15936 17332
rect 2648 17292 15936 17320
rect 2648 17280 2654 17292
rect 15930 17280 15936 17292
rect 15988 17280 15994 17332
rect 16206 17280 16212 17332
rect 16264 17280 16270 17332
rect 1578 17144 1584 17196
rect 1636 17184 1642 17196
rect 2038 17184 2044 17196
rect 1636 17156 2044 17184
rect 1636 17144 1642 17156
rect 2038 17144 2044 17156
rect 2096 17184 2102 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 2096 17156 2421 17184
rect 2096 17144 2102 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 5442 17184 5448 17196
rect 3818 17156 5448 17184
rect 2409 17147 2467 17153
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 6181 17187 6239 17193
rect 6181 17153 6193 17187
rect 6227 17184 6239 17187
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 6227 17156 10425 17184
rect 6227 17153 6239 17156
rect 6181 17147 6239 17153
rect 10413 17153 10425 17156
rect 10459 17153 10471 17187
rect 10413 17147 10471 17153
rect 10686 17144 10692 17196
rect 10744 17144 10750 17196
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11195 17156 11560 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 2682 17076 2688 17128
rect 2740 17076 2746 17128
rect 11532 17125 11560 17156
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 11517 17119 11575 17125
rect 11517 17085 11529 17119
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 4157 16983 4215 16989
rect 4157 16980 4169 16983
rect 4120 16952 4169 16980
rect 4120 16940 4126 16952
rect 4157 16949 4169 16952
rect 4203 16949 4215 16983
rect 4157 16943 4215 16949
rect 5534 16940 5540 16992
rect 5592 16940 5598 16992
rect 11238 16940 11244 16992
rect 11296 16940 11302 16992
rect 11532 16980 11560 17079
rect 11790 17076 11796 17128
rect 11848 17076 11854 17128
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 11940 17088 12848 17116
rect 11940 17076 11946 17088
rect 12820 17048 12848 17088
rect 13354 17076 13360 17128
rect 13412 17076 13418 17128
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 12820 17020 13737 17048
rect 13725 17017 13737 17020
rect 13771 17048 13783 17051
rect 16224 17048 16252 17280
rect 13771 17020 16252 17048
rect 13771 17017 13783 17020
rect 13725 17011 13783 17017
rect 12526 16980 12532 16992
rect 11532 16952 12532 16980
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 13262 16940 13268 16992
rect 13320 16940 13326 16992
rect 13814 16940 13820 16992
rect 13872 16940 13878 16992
rect 1104 16890 17112 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 10214 16890
rect 10266 16838 10278 16890
rect 10330 16838 10342 16890
rect 10394 16838 10406 16890
rect 10458 16838 10470 16890
rect 10522 16838 16214 16890
rect 16266 16838 16278 16890
rect 16330 16838 16342 16890
rect 16394 16838 16406 16890
rect 16458 16838 16470 16890
rect 16522 16838 17112 16890
rect 1104 16816 17112 16838
rect 2777 16779 2835 16785
rect 2777 16745 2789 16779
rect 2823 16776 2835 16779
rect 2866 16776 2872 16788
rect 2823 16748 2872 16776
rect 2823 16745 2835 16748
rect 2777 16739 2835 16745
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 11238 16736 11244 16788
rect 11296 16736 11302 16788
rect 11333 16779 11391 16785
rect 11333 16745 11345 16779
rect 11379 16776 11391 16779
rect 11790 16776 11796 16788
rect 11379 16748 11796 16776
rect 11379 16745 11391 16748
rect 11333 16739 11391 16745
rect 11790 16736 11796 16748
rect 11848 16736 11854 16788
rect 13262 16736 13268 16788
rect 13320 16736 13326 16788
rect 2590 16668 2596 16720
rect 2648 16668 2654 16720
rect 4062 16600 4068 16652
rect 4120 16600 4126 16652
rect 11256 16640 11284 16736
rect 11701 16643 11759 16649
rect 11701 16640 11713 16643
rect 11256 16612 11713 16640
rect 11701 16609 11713 16612
rect 11747 16609 11759 16643
rect 11701 16603 11759 16609
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16640 12035 16643
rect 13280 16640 13308 16736
rect 12023 16612 13308 16640
rect 12023 16609 12035 16612
rect 11977 16603 12035 16609
rect 2130 16532 2136 16584
rect 2188 16572 2194 16584
rect 2869 16575 2927 16581
rect 2869 16572 2881 16575
rect 2188 16544 2881 16572
rect 2188 16532 2194 16544
rect 2869 16541 2881 16544
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3789 16575 3847 16581
rect 3789 16572 3801 16575
rect 3007 16544 3801 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3789 16541 3801 16544
rect 3835 16541 3847 16575
rect 3789 16535 3847 16541
rect 5534 16532 5540 16584
rect 5592 16572 5598 16584
rect 5629 16575 5687 16581
rect 5629 16572 5641 16575
rect 5592 16544 5641 16572
rect 5592 16532 5598 16544
rect 5629 16541 5641 16544
rect 5675 16541 5687 16575
rect 5629 16535 5687 16541
rect 11333 16575 11391 16581
rect 11333 16541 11345 16575
rect 11379 16572 11391 16575
rect 11422 16572 11428 16584
rect 11379 16544 11428 16572
rect 11379 16541 11391 16544
rect 11333 16535 11391 16541
rect 11422 16532 11428 16544
rect 11480 16532 11486 16584
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16541 11575 16575
rect 11517 16535 11575 16541
rect 13725 16575 13783 16581
rect 13725 16541 13737 16575
rect 13771 16572 13783 16575
rect 13814 16572 13820 16584
rect 13771 16544 13820 16572
rect 13771 16541 13783 16544
rect 13725 16535 13783 16541
rect 2314 16464 2320 16516
rect 2372 16464 2378 16516
rect 5442 16504 5448 16516
rect 5290 16476 5448 16504
rect 5442 16464 5448 16476
rect 5500 16464 5506 16516
rect 5534 16396 5540 16448
rect 5592 16396 5598 16448
rect 5810 16396 5816 16448
rect 5868 16396 5874 16448
rect 11532 16436 11560 16535
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 14182 16532 14188 16584
rect 14240 16532 14246 16584
rect 13262 16504 13268 16516
rect 13202 16476 13268 16504
rect 13262 16464 13268 16476
rect 13320 16504 13326 16516
rect 14550 16504 14556 16516
rect 13320 16476 14556 16504
rect 13320 16464 13326 16476
rect 14550 16464 14556 16476
rect 14608 16464 14614 16516
rect 12618 16436 12624 16448
rect 11532 16408 12624 16436
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 12710 16396 12716 16448
rect 12768 16436 12774 16448
rect 13354 16436 13360 16448
rect 12768 16408 13360 16436
rect 12768 16396 12774 16408
rect 13354 16396 13360 16408
rect 13412 16436 13418 16448
rect 13449 16439 13507 16445
rect 13449 16436 13461 16439
rect 13412 16408 13461 16436
rect 13412 16396 13418 16408
rect 13449 16405 13461 16408
rect 13495 16405 13507 16439
rect 13449 16399 13507 16405
rect 13538 16396 13544 16448
rect 13596 16396 13602 16448
rect 14274 16396 14280 16448
rect 14332 16396 14338 16448
rect 1104 16346 17112 16368
rect 1104 16294 7214 16346
rect 7266 16294 7278 16346
rect 7330 16294 7342 16346
rect 7394 16294 7406 16346
rect 7458 16294 7470 16346
rect 7522 16294 13214 16346
rect 13266 16294 13278 16346
rect 13330 16294 13342 16346
rect 13394 16294 13406 16346
rect 13458 16294 13470 16346
rect 13522 16294 17112 16346
rect 1104 16272 17112 16294
rect 2222 16192 2228 16244
rect 2280 16232 2286 16244
rect 5534 16232 5540 16244
rect 2280 16204 5540 16232
rect 2280 16192 2286 16204
rect 1872 16136 2360 16164
rect 934 16056 940 16108
rect 992 16096 998 16108
rect 1872 16105 1900 16136
rect 2332 16108 2360 16136
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 992 16068 1409 16096
rect 992 16056 998 16068
rect 1397 16065 1409 16068
rect 1443 16065 1455 16099
rect 1397 16059 1455 16065
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 1949 16099 2007 16105
rect 1949 16065 1961 16099
rect 1995 16065 2007 16099
rect 1949 16059 2007 16065
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2130 16096 2136 16108
rect 2087 16068 2136 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 1964 16028 1992 16059
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 2222 16056 2228 16108
rect 2280 16056 2286 16108
rect 2314 16056 2320 16108
rect 2372 16056 2378 16108
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16065 2467 16099
rect 2409 16059 2467 16065
rect 2424 16028 2452 16059
rect 2682 16056 2688 16108
rect 2740 16056 2746 16108
rect 2884 16105 2912 16204
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 12897 16167 12955 16173
rect 12897 16133 12909 16167
rect 12943 16164 12955 16167
rect 12943 16136 13308 16164
rect 12943 16133 12955 16136
rect 12897 16127 12955 16133
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 5810 16056 5816 16108
rect 5868 16096 5874 16108
rect 5905 16099 5963 16105
rect 5905 16096 5917 16099
rect 5868 16068 5917 16096
rect 5868 16056 5874 16068
rect 5905 16065 5917 16068
rect 5951 16065 5963 16099
rect 5905 16059 5963 16065
rect 12618 16056 12624 16108
rect 12676 16056 12682 16108
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 12802 16056 12808 16108
rect 12860 16056 12866 16108
rect 13078 16096 13084 16108
rect 13004 16068 13084 16096
rect 1780 16000 2452 16028
rect 12636 16028 12664 16056
rect 13004 16028 13032 16068
rect 13078 16056 13084 16068
rect 13136 16056 13142 16108
rect 13280 16037 13308 16136
rect 13538 16124 13544 16176
rect 13596 16124 13602 16176
rect 14550 16056 14556 16108
rect 14608 16096 14614 16108
rect 14608 16068 14674 16096
rect 14608 16056 14614 16068
rect 12636 16000 13032 16028
rect 13265 16031 13323 16037
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 1780 15960 1808 16000
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 14182 16028 14188 16040
rect 13311 16000 14188 16028
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 14182 15988 14188 16000
rect 14240 15988 14246 16040
rect 1627 15932 1808 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 1780 15904 1808 15932
rect 2501 15963 2559 15969
rect 2501 15929 2513 15963
rect 2547 15960 2559 15963
rect 2774 15960 2780 15972
rect 2547 15932 2780 15960
rect 2547 15929 2559 15932
rect 2501 15923 2559 15929
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 1670 15852 1676 15904
rect 1728 15852 1734 15904
rect 1762 15852 1768 15904
rect 1820 15852 1826 15904
rect 2682 15852 2688 15904
rect 2740 15852 2746 15904
rect 5258 15852 5264 15904
rect 5316 15852 5322 15904
rect 12526 15852 12532 15904
rect 12584 15852 12590 15904
rect 15013 15895 15071 15901
rect 15013 15861 15025 15895
rect 15059 15892 15071 15895
rect 15470 15892 15476 15904
rect 15059 15864 15476 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 1104 15802 17112 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 10214 15802
rect 10266 15750 10278 15802
rect 10330 15750 10342 15802
rect 10394 15750 10406 15802
rect 10458 15750 10470 15802
rect 10522 15750 16214 15802
rect 16266 15750 16278 15802
rect 16330 15750 16342 15802
rect 16394 15750 16406 15802
rect 16458 15750 16470 15802
rect 16522 15750 17112 15802
rect 1104 15728 17112 15750
rect 5800 15691 5858 15697
rect 5800 15657 5812 15691
rect 5846 15688 5858 15691
rect 8573 15691 8631 15697
rect 8573 15688 8585 15691
rect 5846 15660 8585 15688
rect 5846 15657 5858 15660
rect 5800 15651 5858 15657
rect 8573 15657 8585 15660
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 13078 15648 13084 15700
rect 13136 15648 13142 15700
rect 14274 15648 14280 15700
rect 14332 15688 14338 15700
rect 14332 15660 16160 15688
rect 14332 15648 14338 15660
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 9309 15623 9367 15629
rect 5500 15592 5672 15620
rect 5500 15580 5506 15592
rect 1762 15512 1768 15564
rect 1820 15512 1826 15564
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15552 2099 15555
rect 2682 15552 2688 15564
rect 2087 15524 2688 15552
rect 2087 15521 2099 15524
rect 2041 15515 2099 15521
rect 2682 15512 2688 15524
rect 2740 15512 2746 15564
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15521 5595 15555
rect 5644 15552 5672 15592
rect 9309 15589 9321 15623
rect 9355 15620 9367 15623
rect 11422 15620 11428 15632
rect 9355 15592 11428 15620
rect 9355 15589 9367 15592
rect 9309 15583 9367 15589
rect 9324 15552 9352 15583
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 13096 15620 13124 15648
rect 14369 15623 14427 15629
rect 14369 15620 14381 15623
rect 13096 15592 14381 15620
rect 14369 15589 14381 15592
rect 14415 15589 14427 15623
rect 14369 15583 14427 15589
rect 5644 15524 7052 15552
rect 5537 15515 5595 15521
rect 5350 15444 5356 15496
rect 5408 15484 5414 15496
rect 5445 15487 5503 15493
rect 5445 15484 5457 15487
rect 5408 15456 5457 15484
rect 5408 15444 5414 15456
rect 5445 15453 5457 15456
rect 5491 15453 5503 15487
rect 5445 15447 5503 15453
rect 4154 15416 4160 15428
rect 3266 15388 4160 15416
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 4709 15419 4767 15425
rect 4709 15385 4721 15419
rect 4755 15416 4767 15419
rect 5552 15416 5580 15515
rect 6086 15416 6092 15428
rect 4755 15388 6092 15416
rect 4755 15385 4767 15388
rect 4709 15379 4767 15385
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 7024 15416 7052 15524
rect 8588 15524 9352 15552
rect 9401 15555 9459 15561
rect 8588 15493 8616 15524
rect 9401 15521 9413 15555
rect 9447 15552 9459 15555
rect 9447 15524 9720 15552
rect 9447 15521 9459 15524
rect 9401 15515 9459 15521
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 9030 15484 9036 15496
rect 8803 15456 9036 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 9692 15493 9720 15524
rect 15470 15512 15476 15564
rect 15528 15552 15534 15564
rect 16132 15561 16160 15660
rect 15841 15555 15899 15561
rect 15841 15552 15853 15555
rect 15528 15524 15853 15552
rect 15528 15512 15534 15524
rect 15841 15521 15853 15524
rect 15887 15521 15899 15555
rect 15841 15515 15899 15521
rect 16117 15555 16175 15561
rect 16117 15521 16129 15555
rect 16163 15521 16175 15555
rect 16117 15515 16175 15521
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 8294 15416 8300 15428
rect 7024 15402 8300 15416
rect 7038 15388 8300 15402
rect 8294 15376 8300 15388
rect 8352 15376 8358 15428
rect 8662 15376 8668 15428
rect 8720 15416 8726 15428
rect 8941 15419 8999 15425
rect 8941 15416 8953 15419
rect 8720 15388 8953 15416
rect 8720 15376 8726 15388
rect 8941 15385 8953 15388
rect 8987 15385 8999 15419
rect 9876 15416 9904 15447
rect 10962 15416 10968 15428
rect 9876 15388 10968 15416
rect 8941 15379 8999 15385
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 14366 15376 14372 15428
rect 14424 15416 14430 15428
rect 14550 15416 14556 15428
rect 14424 15388 14556 15416
rect 14424 15376 14430 15388
rect 14550 15376 14556 15388
rect 14608 15416 14614 15428
rect 14608 15388 14674 15416
rect 14608 15376 14614 15388
rect 3326 15308 3332 15360
rect 3384 15348 3390 15360
rect 3513 15351 3571 15357
rect 3513 15348 3525 15351
rect 3384 15320 3525 15348
rect 3384 15308 3390 15320
rect 3513 15317 3525 15320
rect 3559 15317 3571 15351
rect 3513 15311 3571 15317
rect 4798 15308 4804 15360
rect 4856 15308 4862 15360
rect 7098 15308 7104 15360
rect 7156 15348 7162 15360
rect 7285 15351 7343 15357
rect 7285 15348 7297 15351
rect 7156 15320 7297 15348
rect 7156 15308 7162 15320
rect 7285 15317 7297 15320
rect 7331 15317 7343 15351
rect 7285 15311 7343 15317
rect 8478 15308 8484 15360
rect 8536 15308 8542 15360
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 9493 15351 9551 15357
rect 9493 15348 9505 15351
rect 9364 15320 9505 15348
rect 9364 15308 9370 15320
rect 9493 15317 9505 15320
rect 9539 15317 9551 15351
rect 9493 15311 9551 15317
rect 9953 15351 10011 15357
rect 9953 15317 9965 15351
rect 9999 15348 10011 15351
rect 11330 15348 11336 15360
rect 9999 15320 11336 15348
rect 9999 15317 10011 15320
rect 9953 15311 10011 15317
rect 11330 15308 11336 15320
rect 11388 15308 11394 15360
rect 11422 15308 11428 15360
rect 11480 15308 11486 15360
rect 1104 15258 17112 15280
rect 1104 15206 7214 15258
rect 7266 15206 7278 15258
rect 7330 15206 7342 15258
rect 7394 15206 7406 15258
rect 7458 15206 7470 15258
rect 7522 15206 13214 15258
rect 13266 15206 13278 15258
rect 13330 15206 13342 15258
rect 13394 15206 13406 15258
rect 13458 15206 13470 15258
rect 13522 15206 17112 15258
rect 1104 15184 17112 15206
rect 5350 15104 5356 15156
rect 5408 15104 5414 15156
rect 8662 15104 8668 15156
rect 8720 15104 8726 15156
rect 9030 15104 9036 15156
rect 9088 15144 9094 15156
rect 9585 15147 9643 15153
rect 9585 15144 9597 15147
rect 9088 15116 9597 15144
rect 9088 15104 9094 15116
rect 9585 15113 9597 15116
rect 9631 15113 9643 15147
rect 9585 15107 9643 15113
rect 10686 15104 10692 15156
rect 10744 15104 10750 15156
rect 13249 15147 13307 15153
rect 13249 15113 13261 15147
rect 13295 15144 13307 15147
rect 13295 15116 13860 15144
rect 13295 15113 13307 15116
rect 13249 15107 13307 15113
rect 1762 15036 1768 15088
rect 1820 15076 1826 15088
rect 2225 15079 2283 15085
rect 2225 15076 2237 15079
rect 1820 15048 2237 15076
rect 1820 15036 1826 15048
rect 2225 15045 2237 15048
rect 2271 15045 2283 15079
rect 2225 15039 2283 15045
rect 3053 15079 3111 15085
rect 3053 15045 3065 15079
rect 3099 15076 3111 15079
rect 3326 15076 3332 15088
rect 3099 15048 3332 15076
rect 3099 15045 3111 15048
rect 3053 15039 3111 15045
rect 3326 15036 3332 15048
rect 3384 15036 3390 15088
rect 7098 15036 7104 15088
rect 7156 15076 7162 15088
rect 7193 15079 7251 15085
rect 7193 15076 7205 15079
rect 7156 15048 7205 15076
rect 7156 15036 7162 15048
rect 7193 15045 7205 15048
rect 7239 15045 7251 15079
rect 7193 15039 7251 15045
rect 8478 15036 8484 15088
rect 8536 15076 8542 15088
rect 9125 15079 9183 15085
rect 9125 15076 9137 15079
rect 8536 15048 9137 15076
rect 8536 15036 8542 15048
rect 9125 15045 9137 15048
rect 9171 15076 9183 15079
rect 10704 15076 10732 15104
rect 13832 15088 13860 15116
rect 14182 15104 14188 15156
rect 14240 15104 14246 15156
rect 9171 15048 9628 15076
rect 10626 15048 10732 15076
rect 9171 15045 9183 15048
rect 9125 15039 9183 15045
rect 9600 15020 9628 15048
rect 10962 15036 10968 15088
rect 11020 15076 11026 15088
rect 13449 15079 13507 15085
rect 13449 15076 13461 15079
rect 11020 15048 13461 15076
rect 11020 15036 11026 15048
rect 13449 15045 13461 15048
rect 13495 15076 13507 15079
rect 13633 15079 13691 15085
rect 13633 15076 13645 15079
rect 13495 15048 13645 15076
rect 13495 15045 13507 15048
rect 13449 15039 13507 15045
rect 13633 15045 13645 15048
rect 13679 15045 13691 15079
rect 13633 15039 13691 15045
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 14200 15076 14228 15104
rect 13872 15048 14228 15076
rect 13872 15036 13878 15048
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 14977 2007 15011
rect 1949 14971 2007 14977
rect 1964 14940 1992 14971
rect 2130 14968 2136 15020
rect 2188 14968 2194 15020
rect 2314 14968 2320 15020
rect 2372 14968 2378 15020
rect 2774 14968 2780 15020
rect 2832 14968 2838 15020
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 4614 15008 4620 15020
rect 4212 14980 4620 15008
rect 4212 14968 4218 14980
rect 4614 14968 4620 14980
rect 4672 14968 4678 15020
rect 4798 14968 4804 15020
rect 4856 14968 4862 15020
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 5353 15011 5411 15017
rect 5353 15008 5365 15011
rect 5316 14980 5365 15008
rect 5316 14968 5322 14980
rect 5353 14977 5365 14980
rect 5399 14977 5411 15011
rect 5353 14971 5411 14977
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 6181 15011 6239 15017
rect 6181 15008 6193 15011
rect 6144 14980 6193 15008
rect 6144 14968 6150 14980
rect 6181 14977 6193 14980
rect 6227 15008 6239 15011
rect 6641 15011 6699 15017
rect 6641 15008 6653 15011
rect 6227 14980 6653 15008
rect 6227 14977 6239 14980
rect 6181 14971 6239 14977
rect 6641 14977 6653 14980
rect 6687 15008 6699 15011
rect 6822 15008 6828 15020
rect 6687 14980 6828 15008
rect 6687 14977 6699 14980
rect 6641 14971 6699 14977
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 8294 14968 8300 15020
rect 8352 14968 8358 15020
rect 8662 14968 8668 15020
rect 8720 14968 8726 15020
rect 8849 15011 8907 15017
rect 8849 14977 8861 15011
rect 8895 15008 8907 15011
rect 8938 15008 8944 15020
rect 8895 14980 8944 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 8938 14968 8944 14980
rect 8996 14968 9002 15020
rect 9030 14968 9036 15020
rect 9088 14968 9094 15020
rect 9222 15011 9280 15017
rect 9222 15008 9234 15011
rect 9140 14980 9234 15008
rect 2222 14940 2228 14952
rect 1964 14912 2228 14940
rect 2222 14900 2228 14912
rect 2280 14900 2286 14952
rect 2332 14940 2360 14968
rect 4525 14943 4583 14949
rect 4525 14940 4537 14943
rect 2332 14912 4537 14940
rect 4525 14909 4537 14912
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 6733 14943 6791 14949
rect 6733 14909 6745 14943
rect 6779 14940 6791 14943
rect 6917 14943 6975 14949
rect 6917 14940 6929 14943
rect 6779 14912 6929 14940
rect 6779 14909 6791 14912
rect 6733 14903 6791 14909
rect 6917 14909 6929 14912
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 8312 14872 8340 14968
rect 8680 14940 8708 14968
rect 9140 14940 9168 14980
rect 9222 14977 9234 14980
rect 9268 14977 9280 15011
rect 9222 14971 9280 14977
rect 9582 14968 9588 15020
rect 9640 14968 9646 15020
rect 11422 14968 11428 15020
rect 11480 15008 11486 15020
rect 11517 15011 11575 15017
rect 11517 15008 11529 15011
rect 11480 14980 11529 15008
rect 11480 14968 11486 14980
rect 11517 14977 11529 14980
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 11773 15011 11831 15017
rect 11773 15008 11785 15011
rect 11664 14980 11785 15008
rect 11664 14968 11670 14980
rect 11773 14977 11785 14980
rect 11819 14977 11831 15011
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 11773 14971 11831 14977
rect 13280 14980 13553 15008
rect 8680 14912 9168 14940
rect 11054 14900 11060 14952
rect 11112 14900 11118 14952
rect 11330 14900 11336 14952
rect 11388 14900 11394 14952
rect 9674 14872 9680 14884
rect 8312 14844 9680 14872
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 13280 14872 13308 14980
rect 13541 14977 13553 14980
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 15008 15439 15011
rect 15930 15008 15936 15020
rect 15427 14980 15936 15008
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 15286 14900 15292 14952
rect 15344 14900 15350 14952
rect 12912 14844 13308 14872
rect 2498 14764 2504 14816
rect 2556 14764 2562 14816
rect 4798 14764 4804 14816
rect 4856 14764 4862 14816
rect 9398 14764 9404 14816
rect 9456 14764 9462 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12802 14804 12808 14816
rect 12492 14776 12808 14804
rect 12492 14764 12498 14776
rect 12802 14764 12808 14776
rect 12860 14804 12866 14816
rect 12912 14813 12940 14844
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12860 14776 12909 14804
rect 12860 14764 12866 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 13280 14813 13308 14844
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 13044 14776 13093 14804
rect 13044 14764 13050 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13081 14767 13139 14773
rect 13265 14807 13323 14813
rect 13265 14773 13277 14807
rect 13311 14773 13323 14807
rect 13265 14767 13323 14773
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 13817 14807 13875 14813
rect 13817 14804 13829 14807
rect 13596 14776 13829 14804
rect 13596 14764 13602 14776
rect 13817 14773 13829 14776
rect 13863 14773 13875 14807
rect 13817 14767 13875 14773
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 15657 14807 15715 14813
rect 15657 14804 15669 14807
rect 15620 14776 15669 14804
rect 15620 14764 15626 14776
rect 15657 14773 15669 14776
rect 15703 14773 15715 14807
rect 15657 14767 15715 14773
rect 1104 14714 17112 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 10214 14714
rect 10266 14662 10278 14714
rect 10330 14662 10342 14714
rect 10394 14662 10406 14714
rect 10458 14662 10470 14714
rect 10522 14662 16214 14714
rect 16266 14662 16278 14714
rect 16330 14662 16342 14714
rect 16394 14662 16406 14714
rect 16458 14662 16470 14714
rect 16522 14662 17112 14714
rect 1104 14640 17112 14662
rect 4798 14560 4804 14612
rect 4856 14560 4862 14612
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 6880 14572 7021 14600
rect 6880 14560 6886 14572
rect 7009 14569 7021 14572
rect 7055 14600 7067 14603
rect 8478 14600 8484 14612
rect 7055 14572 8484 14600
rect 7055 14569 7067 14572
rect 7009 14563 7067 14569
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14396 4675 14399
rect 4816 14396 4844 14560
rect 7116 14473 7144 14572
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14600 10747 14603
rect 11054 14600 11060 14612
rect 10735 14572 11060 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 12250 14600 12256 14612
rect 11480 14572 12256 14600
rect 11480 14560 11486 14572
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 13814 14560 13820 14612
rect 13872 14560 13878 14612
rect 15930 14560 15936 14612
rect 15988 14600 15994 14612
rect 15988 14572 16574 14600
rect 15988 14560 15994 14572
rect 12434 14532 12440 14544
rect 12360 14504 12440 14532
rect 7101 14467 7159 14473
rect 7101 14433 7113 14467
rect 7147 14433 7159 14467
rect 7101 14427 7159 14433
rect 9217 14467 9275 14473
rect 9217 14433 9229 14467
rect 9263 14464 9275 14467
rect 9306 14464 9312 14476
rect 9263 14436 9312 14464
rect 9263 14433 9275 14436
rect 9217 14427 9275 14433
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 11149 14467 11207 14473
rect 11149 14433 11161 14467
rect 11195 14433 11207 14467
rect 11149 14427 11207 14433
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14464 11483 14467
rect 11606 14464 11612 14476
rect 11471 14436 11612 14464
rect 11471 14433 11483 14436
rect 11425 14427 11483 14433
rect 4663 14368 4844 14396
rect 4663 14365 4675 14368
rect 4617 14359 4675 14365
rect 8938 14356 8944 14408
rect 8996 14356 9002 14408
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 11020 14368 11069 14396
rect 11020 14356 11026 14368
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11164 14396 11192 14427
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 12360 14464 12388 14504
rect 12434 14492 12440 14504
rect 12492 14492 12498 14544
rect 16546 14532 16574 14572
rect 16669 14535 16727 14541
rect 16669 14532 16681 14535
rect 16546 14504 16681 14532
rect 16669 14501 16681 14504
rect 16715 14501 16727 14535
rect 16669 14495 16727 14501
rect 12176 14436 12388 14464
rect 12176 14396 12204 14436
rect 11164 14368 12204 14396
rect 11057 14359 11115 14365
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 15562 14405 15568 14408
rect 12437 14399 12495 14405
rect 12437 14396 12449 14399
rect 12308 14368 12449 14396
rect 12308 14356 12314 14368
rect 12437 14365 12449 14368
rect 12483 14365 12495 14399
rect 15289 14399 15347 14405
rect 15289 14396 15301 14399
rect 12437 14359 12495 14365
rect 15120 14368 15301 14396
rect 7368 14331 7426 14337
rect 7368 14297 7380 14331
rect 7414 14328 7426 14331
rect 7834 14328 7840 14340
rect 7414 14300 7840 14328
rect 7414 14297 7426 14300
rect 7368 14291 7426 14297
rect 7834 14288 7840 14300
rect 7892 14288 7898 14340
rect 3970 14220 3976 14272
rect 4028 14220 4034 14272
rect 8481 14263 8539 14269
rect 8481 14229 8493 14263
rect 8527 14260 8539 14263
rect 8956 14260 8984 14356
rect 10686 14328 10692 14340
rect 10442 14300 10692 14328
rect 10686 14288 10692 14300
rect 10744 14288 10750 14340
rect 10980 14260 11008 14356
rect 12704 14331 12762 14337
rect 12704 14297 12716 14331
rect 12750 14328 12762 14331
rect 13078 14328 13084 14340
rect 12750 14300 13084 14328
rect 12750 14297 12762 14300
rect 12704 14291 12762 14297
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 8527 14232 11008 14260
rect 8527 14229 8539 14232
rect 8481 14223 8539 14229
rect 14274 14220 14280 14272
rect 14332 14260 14338 14272
rect 15120 14269 15148 14368
rect 15289 14365 15301 14368
rect 15335 14365 15347 14399
rect 15556 14396 15568 14405
rect 15523 14368 15568 14396
rect 15289 14359 15347 14365
rect 15556 14359 15568 14368
rect 15562 14356 15568 14359
rect 15620 14356 15626 14408
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 14332 14232 15117 14260
rect 14332 14220 14338 14232
rect 15105 14229 15117 14232
rect 15151 14229 15163 14263
rect 15105 14223 15163 14229
rect 1104 14170 17112 14192
rect 1104 14118 7214 14170
rect 7266 14118 7278 14170
rect 7330 14118 7342 14170
rect 7394 14118 7406 14170
rect 7458 14118 7470 14170
rect 7522 14118 13214 14170
rect 13266 14118 13278 14170
rect 13330 14118 13342 14170
rect 13394 14118 13406 14170
rect 13458 14118 13470 14170
rect 13522 14118 17112 14170
rect 1104 14096 17112 14118
rect 3970 14016 3976 14068
rect 4028 14056 4034 14068
rect 4028 14028 4200 14056
rect 4028 14016 4034 14028
rect 4172 13929 4200 14028
rect 7834 14016 7840 14068
rect 7892 14016 7898 14068
rect 8938 14016 8944 14068
rect 8996 14016 9002 14068
rect 13078 14016 13084 14068
rect 13136 14016 13142 14068
rect 13538 14016 13544 14068
rect 13596 14016 13602 14068
rect 15381 14059 15439 14065
rect 15381 14025 15393 14059
rect 15427 14056 15439 14059
rect 15470 14056 15476 14068
rect 15427 14028 15476 14056
rect 15427 14025 15439 14028
rect 15381 14019 15439 14025
rect 15470 14016 15476 14028
rect 15528 14056 15534 14068
rect 15528 14028 15792 14056
rect 15528 14016 15534 14028
rect 4065 13923 4123 13929
rect 4065 13889 4077 13923
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13920 7987 13923
rect 8956 13920 8984 14016
rect 9398 13948 9404 14000
rect 9456 13988 9462 14000
rect 9456 13960 10088 13988
rect 9456 13948 9462 13960
rect 10060 13929 10088 13960
rect 7975 13892 8984 13920
rect 10045 13923 10103 13929
rect 7975 13889 7987 13892
rect 7929 13883 7987 13889
rect 10045 13889 10057 13923
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 4080 13852 4108 13883
rect 12986 13880 12992 13932
rect 13044 13880 13050 13932
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13556 13920 13584 14016
rect 15764 13997 15792 14028
rect 15749 13991 15807 13997
rect 15749 13957 15761 13991
rect 15795 13957 15807 13991
rect 15749 13951 15807 13957
rect 13219 13892 13584 13920
rect 14268 13923 14326 13929
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 14268 13889 14280 13923
rect 14314 13920 14326 13923
rect 14642 13920 14648 13932
rect 14314 13892 14648 13920
rect 14314 13889 14326 13892
rect 14268 13883 14326 13889
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16022 13920 16028 13932
rect 15979 13892 16028 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16022 13880 16028 13892
rect 16080 13880 16086 13932
rect 4433 13855 4491 13861
rect 4433 13852 4445 13855
rect 4080 13824 4445 13852
rect 4433 13821 4445 13824
rect 4479 13821 4491 13855
rect 4433 13815 4491 13821
rect 10134 13812 10140 13864
rect 10192 13812 10198 13864
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 12308 13824 14013 13852
rect 12308 13812 12314 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 3418 13676 3424 13728
rect 3476 13676 3482 13728
rect 13909 13719 13967 13725
rect 13909 13685 13921 13719
rect 13955 13716 13967 13719
rect 14016 13716 14044 13815
rect 14274 13716 14280 13728
rect 13955 13688 14280 13716
rect 13955 13685 13967 13688
rect 13909 13679 13967 13685
rect 14274 13676 14280 13688
rect 14332 13676 14338 13728
rect 15562 13676 15568 13728
rect 15620 13676 15626 13728
rect 1104 13626 17112 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 10214 13626
rect 10266 13574 10278 13626
rect 10330 13574 10342 13626
rect 10394 13574 10406 13626
rect 10458 13574 10470 13626
rect 10522 13574 16214 13626
rect 16266 13574 16278 13626
rect 16330 13574 16342 13626
rect 16394 13574 16406 13626
rect 16458 13574 16470 13626
rect 16522 13574 17112 13626
rect 1104 13552 17112 13574
rect 14642 13472 14648 13524
rect 14700 13472 14706 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15565 13515 15623 13521
rect 15565 13512 15577 13515
rect 15344 13484 15577 13512
rect 15344 13472 15350 13484
rect 9125 13379 9183 13385
rect 9125 13345 9137 13379
rect 9171 13376 9183 13379
rect 9398 13376 9404 13388
rect 9171 13348 9404 13376
rect 9171 13345 9183 13348
rect 9125 13339 9183 13345
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 10410 13336 10416 13388
rect 10468 13376 10474 13388
rect 15396 13385 15424 13484
rect 15565 13481 15577 13484
rect 15611 13481 15623 13515
rect 15565 13475 15623 13481
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 10468 13348 12081 13376
rect 10468 13336 10474 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 3418 13268 3424 13320
rect 3476 13268 3482 13320
rect 6270 13268 6276 13320
rect 6328 13268 6334 13320
rect 10686 13308 10692 13320
rect 10534 13280 10692 13308
rect 10686 13268 10692 13280
rect 10744 13308 10750 13320
rect 12434 13308 12440 13320
rect 10744 13280 12440 13308
rect 10744 13268 10750 13280
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 13814 13268 13820 13320
rect 13872 13268 13878 13320
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14875 13280 15025 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 15013 13277 15025 13280
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 15197 13311 15255 13317
rect 15197 13277 15209 13311
rect 15243 13277 15255 13311
rect 15197 13271 15255 13277
rect 6546 13200 6552 13252
rect 6604 13200 6610 13252
rect 8294 13240 8300 13252
rect 6932 13212 7038 13240
rect 7944 13212 8300 13240
rect 3418 13132 3424 13184
rect 3476 13132 3482 13184
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 6932 13172 6960 13212
rect 7944 13172 7972 13212
rect 8294 13200 8300 13212
rect 8352 13240 8358 13252
rect 8846 13240 8852 13252
rect 8352 13212 8852 13240
rect 8352 13200 8358 13212
rect 8846 13200 8852 13212
rect 8904 13200 8910 13252
rect 9306 13200 9312 13252
rect 9364 13240 9370 13252
rect 9401 13243 9459 13249
rect 9401 13240 9413 13243
rect 9364 13212 9413 13240
rect 9364 13200 9370 13212
rect 9401 13209 9413 13212
rect 9447 13209 9459 13243
rect 9401 13203 9459 13209
rect 13538 13200 13544 13252
rect 13596 13200 13602 13252
rect 15212 13240 15240 13271
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 15562 13268 15568 13320
rect 15620 13268 15626 13320
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13308 15715 13311
rect 15703 13280 16068 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 15580 13240 15608 13268
rect 15212 13212 15608 13240
rect 16040 13184 16068 13280
rect 4672 13144 7972 13172
rect 4672 13132 4678 13144
rect 8018 13132 8024 13184
rect 8076 13132 8082 13184
rect 10870 13132 10876 13184
rect 10928 13132 10934 13184
rect 16022 13132 16028 13184
rect 16080 13132 16086 13184
rect 1104 13082 17112 13104
rect 1104 13030 7214 13082
rect 7266 13030 7278 13082
rect 7330 13030 7342 13082
rect 7394 13030 7406 13082
rect 7458 13030 7470 13082
rect 7522 13030 13214 13082
rect 13266 13030 13278 13082
rect 13330 13030 13342 13082
rect 13394 13030 13406 13082
rect 13458 13030 13470 13082
rect 13522 13030 17112 13082
rect 1104 13008 17112 13030
rect 7193 12971 7251 12977
rect 7193 12937 7205 12971
rect 7239 12968 7251 12971
rect 8018 12968 8024 12980
rect 7239 12940 7420 12968
rect 7239 12937 7251 12940
rect 7193 12931 7251 12937
rect 2498 12860 2504 12912
rect 2556 12900 2562 12912
rect 2685 12903 2743 12909
rect 2685 12900 2697 12903
rect 2556 12872 2697 12900
rect 2556 12860 2562 12872
rect 2685 12869 2697 12872
rect 2731 12869 2743 12903
rect 2685 12863 2743 12869
rect 5000 12872 7052 12900
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 2915 12804 3157 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3145 12801 3157 12804
rect 3191 12832 3203 12835
rect 4890 12832 4896 12844
rect 3191 12804 4896 12832
rect 3191 12801 3203 12804
rect 3145 12795 3203 12801
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 5000 12841 5028 12872
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12801 5043 12835
rect 4985 12795 5043 12801
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 6270 12832 6276 12844
rect 5675 12804 6276 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 5718 12724 5724 12776
rect 5776 12724 5782 12776
rect 6914 12724 6920 12776
rect 6972 12724 6978 12776
rect 7024 12764 7052 12872
rect 7098 12792 7104 12844
rect 7156 12792 7162 12844
rect 7392 12841 7420 12940
rect 7668 12940 8024 12968
rect 7668 12909 7696 12940
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 9306 12928 9312 12980
rect 9364 12928 9370 12980
rect 10594 12968 10600 12980
rect 9876 12940 10600 12968
rect 7653 12903 7711 12909
rect 7653 12869 7665 12903
rect 7699 12869 7711 12903
rect 7653 12863 7711 12869
rect 8294 12860 8300 12912
rect 8352 12860 8358 12912
rect 9876 12900 9904 12940
rect 10594 12928 10600 12940
rect 10652 12928 10658 12980
rect 10689 12971 10747 12977
rect 10689 12937 10701 12971
rect 10735 12968 10747 12971
rect 10778 12968 10784 12980
rect 10735 12940 10784 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 10965 12971 11023 12977
rect 10965 12937 10977 12971
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 13265 12971 13323 12977
rect 13265 12937 13277 12971
rect 13311 12968 13323 12971
rect 13538 12968 13544 12980
rect 13311 12940 13544 12968
rect 13311 12937 13323 12940
rect 13265 12931 13323 12937
rect 9416 12872 9904 12900
rect 9953 12903 10011 12909
rect 9416 12841 9444 12872
rect 9953 12869 9965 12903
rect 9999 12900 10011 12903
rect 10980 12900 11008 12931
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 11793 12903 11851 12909
rect 11793 12900 11805 12903
rect 9999 12872 10916 12900
rect 10980 12872 11805 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 9217 12835 9275 12841
rect 9217 12801 9229 12835
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9232 12764 9260 12795
rect 9490 12792 9496 12844
rect 9548 12832 9554 12844
rect 9717 12835 9775 12841
rect 9717 12832 9729 12835
rect 9548 12804 9729 12832
rect 9548 12792 9554 12804
rect 9717 12801 9729 12804
rect 9763 12801 9775 12835
rect 9717 12795 9775 12801
rect 9858 12792 9864 12844
rect 9916 12792 9922 12844
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 10410 12832 10416 12844
rect 10183 12804 10416 12832
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 7024 12736 8708 12764
rect 9232 12736 9720 12764
rect 5258 12656 5264 12708
rect 5316 12656 5322 12708
rect 5902 12656 5908 12708
rect 5960 12696 5966 12708
rect 6638 12696 6644 12708
rect 5960 12668 6644 12696
rect 5960 12656 5966 12668
rect 6638 12656 6644 12668
rect 6696 12656 6702 12708
rect 8680 12696 8708 12736
rect 9585 12699 9643 12705
rect 8680 12668 9260 12696
rect 3050 12588 3056 12640
rect 3108 12588 3114 12640
rect 4798 12588 4804 12640
rect 4856 12588 4862 12640
rect 6454 12588 6460 12640
rect 6512 12588 6518 12640
rect 9122 12588 9128 12640
rect 9180 12588 9186 12640
rect 9232 12628 9260 12668
rect 9585 12665 9597 12699
rect 9631 12665 9643 12699
rect 9692 12696 9720 12736
rect 10152 12696 10180 12795
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10778 12792 10784 12844
rect 10836 12792 10842 12844
rect 10888 12832 10916 12872
rect 11793 12869 11805 12872
rect 11839 12869 11851 12903
rect 11793 12863 11851 12869
rect 12434 12860 12440 12912
rect 12492 12860 12498 12912
rect 15010 12860 15016 12912
rect 15068 12900 15074 12912
rect 15105 12903 15163 12909
rect 15105 12900 15117 12903
rect 15068 12872 15117 12900
rect 15068 12860 15074 12872
rect 15105 12869 15117 12872
rect 15151 12869 15163 12903
rect 15105 12863 15163 12869
rect 15194 12860 15200 12912
rect 15252 12900 15258 12912
rect 15305 12903 15363 12909
rect 15305 12900 15317 12903
rect 15252 12872 15317 12900
rect 15252 12860 15258 12872
rect 15305 12869 15317 12872
rect 15351 12869 15363 12903
rect 15305 12863 15363 12869
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 10888 12804 11529 12832
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 10229 12767 10287 12773
rect 10229 12733 10241 12767
rect 10275 12733 10287 12767
rect 11532 12764 11560 12795
rect 15838 12792 15844 12844
rect 15896 12832 15902 12844
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 15896 12804 16313 12832
rect 15896 12792 15902 12804
rect 16301 12801 16313 12804
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 12526 12764 12532 12776
rect 11532 12736 12532 12764
rect 10229 12727 10287 12733
rect 9692 12668 10180 12696
rect 9585 12659 9643 12665
rect 9600 12628 9628 12659
rect 9232 12600 9628 12628
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 10244 12628 10272 12727
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 10594 12656 10600 12708
rect 10652 12656 10658 12708
rect 12250 12628 12256 12640
rect 9916 12600 12256 12628
rect 9916 12588 9922 12600
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 14274 12588 14280 12640
rect 14332 12588 14338 12640
rect 15286 12588 15292 12640
rect 15344 12588 15350 12640
rect 15473 12631 15531 12637
rect 15473 12597 15485 12631
rect 15519 12628 15531 12631
rect 16022 12628 16028 12640
rect 15519 12600 16028 12628
rect 15519 12597 15531 12600
rect 15473 12591 15531 12597
rect 16022 12588 16028 12600
rect 16080 12588 16086 12640
rect 16114 12588 16120 12640
rect 16172 12628 16178 12640
rect 16485 12631 16543 12637
rect 16485 12628 16497 12631
rect 16172 12600 16497 12628
rect 16172 12588 16178 12600
rect 16485 12597 16497 12600
rect 16531 12597 16543 12631
rect 16485 12591 16543 12597
rect 1104 12538 17112 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 10214 12538
rect 10266 12486 10278 12538
rect 10330 12486 10342 12538
rect 10394 12486 10406 12538
rect 10458 12486 10470 12538
rect 10522 12486 16214 12538
rect 16266 12486 16278 12538
rect 16330 12486 16342 12538
rect 16394 12486 16406 12538
rect 16458 12486 16470 12538
rect 16522 12486 17112 12538
rect 1104 12464 17112 12486
rect 6546 12384 6552 12436
rect 6604 12424 6610 12436
rect 6641 12427 6699 12433
rect 6641 12424 6653 12427
rect 6604 12396 6653 12424
rect 6604 12384 6610 12396
rect 6641 12393 6653 12396
rect 6687 12393 6699 12427
rect 6641 12387 6699 12393
rect 12250 12384 12256 12436
rect 12308 12384 12314 12436
rect 12437 12427 12495 12433
rect 12437 12393 12449 12427
rect 12483 12424 12495 12427
rect 13814 12424 13820 12436
rect 12483 12396 13820 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 14415 12396 16068 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 6089 12359 6147 12365
rect 6089 12325 6101 12359
rect 6135 12356 6147 12359
rect 6270 12356 6276 12368
rect 6135 12328 6276 12356
rect 6135 12325 6147 12328
rect 6089 12319 6147 12325
rect 6270 12316 6276 12328
rect 6328 12356 6334 12368
rect 7098 12356 7104 12368
rect 6328 12328 7104 12356
rect 6328 12316 6334 12328
rect 7098 12316 7104 12328
rect 7156 12316 7162 12368
rect 12526 12316 12532 12368
rect 12584 12316 12590 12368
rect 13078 12316 13084 12368
rect 13136 12316 13142 12368
rect 1670 12248 1676 12300
rect 1728 12288 1734 12300
rect 1857 12291 1915 12297
rect 1857 12288 1869 12291
rect 1728 12260 1869 12288
rect 1728 12248 1734 12260
rect 1857 12257 1869 12260
rect 1903 12257 1915 12291
rect 1857 12251 1915 12257
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10505 12291 10563 12297
rect 10505 12288 10517 12291
rect 10192 12260 10517 12288
rect 10192 12248 10198 12260
rect 10505 12257 10517 12260
rect 10551 12257 10563 12291
rect 10505 12251 10563 12257
rect 10778 12248 10784 12300
rect 10836 12248 10842 12300
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 4976 12223 5034 12229
rect 4976 12189 4988 12223
rect 5022 12220 5034 12223
rect 5258 12220 5264 12232
rect 5022 12192 5264 12220
rect 5022 12189 5034 12192
rect 4976 12183 5034 12189
rect 5258 12180 5264 12192
rect 5316 12180 5322 12232
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 12544 12229 12572 12316
rect 13096 12288 13124 12316
rect 14918 12288 14924 12300
rect 13096 12260 13584 12288
rect 13556 12229 13584 12260
rect 14200 12260 14924 12288
rect 14200 12229 14228 12260
rect 14918 12248 14924 12260
rect 14976 12248 14982 12300
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 6512 12192 6837 12220
rect 6512 12180 6518 12192
rect 6825 12189 6837 12192
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12189 12587 12223
rect 13357 12223 13415 12229
rect 13357 12220 13369 12223
rect 12529 12183 12587 12189
rect 12728 12192 13369 12220
rect 2130 12112 2136 12164
rect 2188 12112 2194 12164
rect 3694 12152 3700 12164
rect 3358 12124 3700 12152
rect 3694 12112 3700 12124
rect 3752 12152 3758 12164
rect 4614 12152 4620 12164
rect 3752 12124 4620 12152
rect 3752 12112 3758 12124
rect 4614 12112 4620 12124
rect 4672 12112 4678 12164
rect 12434 12152 12440 12164
rect 12006 12124 12440 12152
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 12728 12096 12756 12192
rect 13357 12189 13369 12192
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12189 13599 12223
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13541 12183 13599 12189
rect 13740 12192 14105 12220
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 3605 12087 3663 12093
rect 3605 12084 3617 12087
rect 3476 12056 3617 12084
rect 3476 12044 3482 12056
rect 3605 12053 3617 12056
rect 3651 12053 3663 12087
rect 3605 12047 3663 12053
rect 12710 12044 12716 12096
rect 12768 12044 12774 12096
rect 13372 12084 13400 12183
rect 13740 12164 13768 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14185 12223 14243 12229
rect 14185 12189 14197 12223
rect 14231 12189 14243 12223
rect 14185 12183 14243 12189
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 16040 12229 16068 12396
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 14332 12192 15945 12220
rect 14332 12180 14338 12192
rect 15933 12189 15945 12192
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16206 12180 16212 12232
rect 16264 12180 16270 12232
rect 13722 12112 13728 12164
rect 13780 12112 13786 12164
rect 14369 12155 14427 12161
rect 14369 12121 14381 12155
rect 14415 12121 14427 12155
rect 14369 12115 14427 12121
rect 14182 12084 14188 12096
rect 13372 12056 14188 12084
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14384 12084 14412 12115
rect 15286 12112 15292 12164
rect 15344 12112 15350 12164
rect 15688 12155 15746 12161
rect 15688 12121 15700 12155
rect 15734 12152 15746 12155
rect 16117 12155 16175 12161
rect 16117 12152 16129 12155
rect 15734 12124 16129 12152
rect 15734 12121 15746 12124
rect 15688 12115 15746 12121
rect 16117 12121 16129 12124
rect 16163 12121 16175 12155
rect 16117 12115 16175 12121
rect 14553 12087 14611 12093
rect 14553 12084 14565 12087
rect 14384 12056 14565 12084
rect 14553 12053 14565 12056
rect 14599 12084 14611 12087
rect 15304 12084 15332 12112
rect 14599 12056 15332 12084
rect 14599 12053 14611 12056
rect 14553 12047 14611 12053
rect 1104 11994 17112 12016
rect 1104 11942 7214 11994
rect 7266 11942 7278 11994
rect 7330 11942 7342 11994
rect 7394 11942 7406 11994
rect 7458 11942 7470 11994
rect 7522 11942 13214 11994
rect 13266 11942 13278 11994
rect 13330 11942 13342 11994
rect 13394 11942 13406 11994
rect 13458 11942 13470 11994
rect 13522 11942 17112 11994
rect 1104 11920 17112 11942
rect 3418 11880 3424 11892
rect 3160 11852 3424 11880
rect 3160 11821 3188 11852
rect 3418 11840 3424 11852
rect 3476 11840 3482 11892
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 5269 11883 5327 11889
rect 5269 11880 5281 11883
rect 4764 11852 5281 11880
rect 4764 11840 4770 11852
rect 5269 11849 5281 11852
rect 5315 11849 5327 11883
rect 5269 11843 5327 11849
rect 6914 11840 6920 11892
rect 6972 11880 6978 11892
rect 13078 11880 13084 11892
rect 6972 11852 7788 11880
rect 6972 11840 6978 11852
rect 3145 11815 3203 11821
rect 3145 11781 3157 11815
rect 3191 11781 3203 11815
rect 4614 11812 4620 11824
rect 4370 11784 4620 11812
rect 3145 11775 3203 11781
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 7098 11772 7104 11824
rect 7156 11812 7162 11824
rect 7561 11815 7619 11821
rect 7561 11812 7573 11815
rect 7156 11784 7573 11812
rect 7156 11772 7162 11784
rect 7561 11781 7573 11784
rect 7607 11781 7619 11815
rect 7561 11775 7619 11781
rect 7760 11812 7788 11852
rect 12912 11852 13084 11880
rect 7760 11784 9260 11812
rect 2866 11704 2872 11756
rect 2924 11704 2930 11756
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 4632 11716 4721 11744
rect 4154 11568 4160 11620
rect 4212 11568 4218 11620
rect 4172 11540 4200 11568
rect 4632 11549 4660 11716
rect 4709 11713 4721 11716
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 4798 11704 4804 11756
rect 4856 11704 4862 11756
rect 4890 11704 4896 11756
rect 4948 11704 4954 11756
rect 4982 11704 4988 11756
rect 5040 11704 5046 11756
rect 5082 11747 5140 11753
rect 5082 11713 5094 11747
rect 5128 11713 5140 11747
rect 5082 11707 5140 11713
rect 4816 11676 4844 11704
rect 5092 11676 5120 11707
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 6696 11716 7021 11744
rect 6696 11704 6702 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7009 11707 7067 11713
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11744 7251 11747
rect 7377 11747 7435 11753
rect 7377 11744 7389 11747
rect 7239 11716 7389 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 7377 11713 7389 11716
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 4816 11648 5120 11676
rect 7392 11676 7420 11707
rect 7650 11704 7656 11756
rect 7708 11704 7714 11756
rect 7760 11753 7788 11784
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 9122 11704 9128 11756
rect 9180 11704 9186 11756
rect 9232 11744 9260 11784
rect 9674 11772 9680 11824
rect 9732 11812 9738 11824
rect 9732 11784 12848 11812
rect 9732 11772 9738 11784
rect 12820 11756 12848 11784
rect 9858 11744 9864 11756
rect 9232 11716 9864 11744
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11744 10931 11747
rect 10919 11716 11192 11744
rect 10919 11713 10931 11716
rect 10873 11707 10931 11713
rect 9140 11676 9168 11704
rect 7392 11648 9168 11676
rect 11164 11620 11192 11716
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 12802 11704 12808 11756
rect 12860 11704 12866 11756
rect 12912 11753 12940 11852
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 14240 11852 14381 11880
rect 14240 11840 14246 11852
rect 14369 11849 14381 11852
rect 14415 11880 14427 11883
rect 15102 11880 15108 11892
rect 14415 11852 15108 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 14274 11812 14280 11824
rect 13004 11784 14280 11812
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 13004 11685 13032 11784
rect 14274 11772 14280 11784
rect 14332 11812 14338 11824
rect 14829 11815 14887 11821
rect 14829 11812 14841 11815
rect 14332 11784 14841 11812
rect 14332 11772 14338 11784
rect 14829 11781 14841 11784
rect 14875 11812 14887 11815
rect 14875 11784 15056 11812
rect 14875 11781 14887 11784
rect 14829 11775 14887 11781
rect 13256 11747 13314 11753
rect 13256 11713 13268 11747
rect 13302 11744 13314 11747
rect 13538 11744 13544 11756
rect 13302 11716 13544 11744
rect 13302 11713 13314 11716
rect 13256 11707 13314 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 15028 11753 15056 11784
rect 15286 11753 15292 11756
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 15280 11707 15292 11753
rect 15286 11704 15292 11707
rect 15344 11704 15350 11756
rect 12989 11679 13047 11685
rect 12989 11676 13001 11679
rect 12544 11648 13001 11676
rect 11146 11568 11152 11620
rect 11204 11568 11210 11620
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4172 11512 4629 11540
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 7006 11500 7012 11552
rect 7064 11500 7070 11552
rect 7926 11500 7932 11552
rect 7984 11500 7990 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 8904 11512 9413 11540
rect 8904 11500 8910 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11540 11023 11543
rect 11330 11540 11336 11552
rect 11011 11512 11336 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 11422 11500 11428 11552
rect 11480 11540 11486 11552
rect 12544 11549 12572 11648
rect 12989 11645 13001 11648
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 12529 11543 12587 11549
rect 12529 11540 12541 11543
rect 11480 11512 12541 11540
rect 11480 11500 11486 11512
rect 12529 11509 12541 11512
rect 12575 11509 12587 11543
rect 12529 11503 12587 11509
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13262 11540 13268 11552
rect 12943 11512 13268 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 15068 11512 16405 11540
rect 15068 11500 15074 11512
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 1104 11450 17112 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 10214 11450
rect 10266 11398 10278 11450
rect 10330 11398 10342 11450
rect 10394 11398 10406 11450
rect 10458 11398 10470 11450
rect 10522 11398 16214 11450
rect 16266 11398 16278 11450
rect 16330 11398 16342 11450
rect 16394 11398 16406 11450
rect 16458 11398 16470 11450
rect 16522 11398 17112 11450
rect 1104 11376 17112 11398
rect 2130 11296 2136 11348
rect 2188 11336 2194 11348
rect 2593 11339 2651 11345
rect 2593 11336 2605 11339
rect 2188 11308 2605 11336
rect 2188 11296 2194 11308
rect 2593 11305 2605 11308
rect 2639 11305 2651 11339
rect 2593 11299 2651 11305
rect 7006 11296 7012 11348
rect 7064 11296 7070 11348
rect 7926 11296 7932 11348
rect 7984 11336 7990 11348
rect 11146 11336 11152 11348
rect 7984 11308 11152 11336
rect 7984 11296 7990 11308
rect 4614 11228 4620 11280
rect 4672 11228 4678 11280
rect 2608 11172 4384 11200
rect 2406 11092 2412 11144
rect 2464 11092 2470 11144
rect 2608 11141 2636 11172
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11101 2651 11135
rect 2593 11095 2651 11101
rect 4062 11092 4068 11144
rect 4120 11092 4126 11144
rect 4356 11076 4384 11172
rect 5718 11160 5724 11212
rect 5776 11200 5782 11212
rect 6181 11203 6239 11209
rect 6181 11200 6193 11203
rect 5776 11172 6193 11200
rect 5776 11160 5782 11172
rect 6181 11169 6193 11172
rect 6227 11200 6239 11203
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 6227 11172 6377 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 6365 11169 6377 11172
rect 6411 11169 6423 11203
rect 7024 11200 7052 11296
rect 9876 11209 9904 11308
rect 11146 11296 11152 11308
rect 11204 11296 11210 11348
rect 11330 11296 11336 11348
rect 11388 11296 11394 11348
rect 13262 11296 13268 11348
rect 13320 11296 13326 11348
rect 13538 11296 13544 11348
rect 13596 11296 13602 11348
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 15344 11308 15485 11336
rect 15344 11296 15350 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 7024 11172 7205 11200
rect 6365 11163 6423 11169
rect 7193 11169 7205 11172
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 9861 11203 9919 11209
rect 9861 11169 9873 11203
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 4485 11135 4543 11141
rect 4485 11101 4497 11135
rect 4531 11132 4543 11135
rect 4798 11132 4804 11144
rect 4531 11104 4804 11132
rect 4531 11101 4543 11104
rect 4485 11095 4543 11101
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 4982 11092 4988 11144
rect 5040 11092 5046 11144
rect 5994 11092 6000 11144
rect 6052 11092 6058 11144
rect 6273 11135 6331 11141
rect 6273 11101 6285 11135
rect 6319 11101 6331 11135
rect 6273 11095 6331 11101
rect 6457 11135 6515 11141
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 6822 11132 6828 11144
rect 6503 11104 6828 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 4249 11067 4307 11073
rect 4249 11033 4261 11067
rect 4295 11033 4307 11067
rect 4249 11027 4307 11033
rect 4264 10996 4292 11027
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 5000 11064 5028 11092
rect 4396 11036 5028 11064
rect 4396 11024 4402 11036
rect 6288 11008 6316 11095
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6880 11104 6929 11132
rect 6880 11092 6886 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 11348 11132 11376 11296
rect 11609 11203 11667 11209
rect 11609 11169 11621 11203
rect 11655 11200 11667 11203
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11655 11172 11989 11200
rect 11655 11169 11667 11172
rect 11609 11163 11667 11169
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 11977 11163 12035 11169
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 12492 11172 13124 11200
rect 12492 11160 12498 11172
rect 13096 11144 13124 11172
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11348 11104 11713 11132
rect 6917 11095 6975 11101
rect 11701 11101 11713 11104
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 13078 11092 13084 11144
rect 13136 11092 13142 11144
rect 13280 11132 13308 11296
rect 15013 11203 15071 11209
rect 15013 11169 15025 11203
rect 15059 11200 15071 11203
rect 15194 11200 15200 11212
rect 15059 11172 15200 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13280 11104 13553 11132
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 15028 11132 15056 11163
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 13780 11104 15056 11132
rect 15105 11135 15163 11141
rect 13780 11092 13786 11104
rect 15105 11101 15117 11135
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 8846 11064 8852 11076
rect 8418 11036 8852 11064
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 10134 11024 10140 11076
rect 10192 11024 10198 11076
rect 12434 11064 12440 11076
rect 11362 11036 12440 11064
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 15010 11024 15016 11076
rect 15068 11064 15074 11076
rect 15120 11064 15148 11095
rect 15068 11036 15148 11064
rect 15068 11024 15074 11036
rect 4706 10996 4712 11008
rect 4264 10968 4712 10996
rect 4706 10956 4712 10968
rect 4764 10996 4770 11008
rect 4890 10996 4896 11008
rect 4764 10968 4896 10996
rect 4764 10956 4770 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5810 10956 5816 11008
rect 5868 10956 5874 11008
rect 6270 10956 6276 11008
rect 6328 10956 6334 11008
rect 8662 10956 8668 11008
rect 8720 10956 8726 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 13449 10999 13507 11005
rect 13449 10996 13461 10999
rect 12676 10968 13461 10996
rect 12676 10956 12682 10968
rect 13449 10965 13461 10968
rect 13495 10965 13507 10999
rect 13449 10959 13507 10965
rect 1104 10906 17112 10928
rect 1104 10854 7214 10906
rect 7266 10854 7278 10906
rect 7330 10854 7342 10906
rect 7394 10854 7406 10906
rect 7458 10854 7470 10906
rect 7522 10854 13214 10906
rect 13266 10854 13278 10906
rect 13330 10854 13342 10906
rect 13394 10854 13406 10906
rect 13458 10854 13470 10906
rect 13522 10854 17112 10906
rect 1104 10832 17112 10854
rect 4338 10792 4344 10804
rect 3068 10764 4344 10792
rect 3068 10733 3096 10764
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 4798 10752 4804 10804
rect 4856 10752 4862 10804
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 6052 10764 6377 10792
rect 6052 10752 6058 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 7650 10752 7656 10804
rect 7708 10752 7714 10804
rect 9858 10752 9864 10804
rect 9916 10752 9922 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 10192 10764 10517 10792
rect 10192 10752 10198 10764
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 10505 10755 10563 10761
rect 3053 10727 3111 10733
rect 3053 10693 3065 10727
rect 3099 10693 3111 10727
rect 4816 10724 4844 10752
rect 3053 10687 3111 10693
rect 4080 10696 4844 10724
rect 6733 10727 6791 10733
rect 2774 10616 2780 10668
rect 2832 10616 2838 10668
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10625 3019 10659
rect 2961 10619 3019 10625
rect 3197 10659 3255 10665
rect 3197 10625 3209 10659
rect 3243 10656 3255 10659
rect 4080 10656 4108 10696
rect 6733 10693 6745 10727
rect 6779 10724 6791 10727
rect 6822 10724 6828 10736
rect 6779 10696 6828 10724
rect 6779 10693 6791 10696
rect 6733 10687 6791 10693
rect 3243 10628 4108 10656
rect 3243 10625 3255 10628
rect 3197 10619 3255 10625
rect 934 10548 940 10600
rect 992 10588 998 10600
rect 1397 10591 1455 10597
rect 1397 10588 1409 10591
rect 992 10560 1409 10588
rect 992 10548 998 10560
rect 1397 10557 1409 10560
rect 1443 10557 1455 10591
rect 2976 10588 3004 10619
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4672 10628 4813 10656
rect 4672 10616 4678 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 5068 10659 5126 10665
rect 5068 10625 5080 10659
rect 5114 10656 5126 10659
rect 5534 10656 5540 10668
rect 5114 10628 5540 10656
rect 5114 10625 5126 10628
rect 5068 10619 5126 10625
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 6270 10616 6276 10668
rect 6328 10656 6334 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6328 10628 6561 10656
rect 6328 10616 6334 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 4706 10588 4712 10600
rect 2976 10560 4712 10588
rect 1397 10551 1455 10557
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 6181 10523 6239 10529
rect 6181 10489 6193 10523
rect 6227 10520 6239 10523
rect 6748 10520 6776 10687
rect 6822 10684 6828 10696
rect 6880 10724 6886 10736
rect 7668 10724 7696 10752
rect 6880 10696 7696 10724
rect 6880 10684 6886 10696
rect 7668 10656 7696 10696
rect 8389 10727 8447 10733
rect 8389 10693 8401 10727
rect 8435 10724 8447 10727
rect 8662 10724 8668 10736
rect 8435 10696 8668 10724
rect 8435 10693 8447 10696
rect 8389 10687 8447 10693
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 8846 10684 8852 10736
rect 8904 10684 8910 10736
rect 12250 10684 12256 10736
rect 12308 10724 12314 10736
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 12308 10696 15025 10724
rect 12308 10684 12314 10696
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7668 10628 7757 10656
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 8113 10591 8171 10597
rect 8113 10588 8125 10591
rect 7883 10560 8125 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 8113 10557 8125 10560
rect 8159 10557 8171 10591
rect 10704 10588 10732 10619
rect 12894 10616 12900 10668
rect 12952 10616 12958 10668
rect 14292 10665 14320 10696
rect 15013 10693 15025 10696
rect 15059 10693 15071 10727
rect 15013 10687 15071 10693
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 14826 10616 14832 10668
rect 14884 10616 14890 10668
rect 15102 10616 15108 10668
rect 15160 10616 15166 10668
rect 15194 10616 15200 10668
rect 15252 10665 15258 10668
rect 15252 10656 15260 10665
rect 15470 10656 15476 10668
rect 15252 10628 15476 10656
rect 15252 10619 15260 10628
rect 15252 10616 15258 10619
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10704 10560 10793 10588
rect 8113 10551 8171 10557
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 11238 10548 11244 10600
rect 11296 10548 11302 10600
rect 13078 10548 13084 10600
rect 13136 10588 13142 10600
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 13136 10560 13185 10588
rect 13136 10548 13142 10560
rect 13173 10557 13185 10560
rect 13219 10588 13231 10591
rect 13998 10588 14004 10600
rect 13219 10560 14004 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 15838 10548 15844 10600
rect 15896 10548 15902 10600
rect 6227 10492 6776 10520
rect 10965 10523 11023 10529
rect 6227 10489 6239 10492
rect 6181 10483 6239 10489
rect 10965 10489 10977 10523
rect 11011 10520 11023 10523
rect 15381 10523 15439 10529
rect 11011 10492 11560 10520
rect 11011 10489 11023 10492
rect 10965 10483 11023 10489
rect 11532 10464 11560 10492
rect 15381 10489 15393 10523
rect 15427 10520 15439 10523
rect 15856 10520 15884 10548
rect 15427 10492 15884 10520
rect 15427 10489 15439 10492
rect 15381 10483 15439 10489
rect 3326 10412 3332 10464
rect 3384 10412 3390 10464
rect 11514 10412 11520 10464
rect 11572 10412 11578 10464
rect 13354 10412 13360 10464
rect 13412 10412 13418 10464
rect 14182 10412 14188 10464
rect 14240 10412 14246 10464
rect 1104 10362 17112 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 10214 10362
rect 10266 10310 10278 10362
rect 10330 10310 10342 10362
rect 10394 10310 10406 10362
rect 10458 10310 10470 10362
rect 10522 10310 16214 10362
rect 16266 10310 16278 10362
rect 16330 10310 16342 10362
rect 16394 10310 16406 10362
rect 16458 10310 16470 10362
rect 16522 10310 17112 10362
rect 1104 10288 17112 10310
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3513 10251 3571 10257
rect 3513 10248 3525 10251
rect 3108 10220 3525 10248
rect 3108 10208 3114 10220
rect 3513 10217 3525 10220
rect 3559 10217 3571 10251
rect 3513 10211 3571 10217
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 12618 10248 12624 10260
rect 11716 10220 12624 10248
rect 2866 10140 2872 10192
rect 2924 10180 2930 10192
rect 2924 10152 3832 10180
rect 2924 10140 2930 10152
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 1627 10084 3648 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 3620 10053 3648 10084
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10013 3663 10047
rect 3804 10044 3832 10152
rect 4614 10140 4620 10192
rect 4672 10140 4678 10192
rect 11238 10180 11244 10192
rect 10796 10152 11244 10180
rect 4062 10044 4068 10056
rect 3804 10016 4068 10044
rect 3605 10007 3663 10013
rect 1854 9936 1860 9988
rect 1912 9936 1918 9988
rect 3620 9976 3648 10007
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4485 10047 4543 10053
rect 4485 10044 4497 10047
rect 4172 10016 4497 10044
rect 4172 9976 4200 10016
rect 4485 10013 4497 10016
rect 4531 10044 4543 10047
rect 4798 10044 4804 10056
rect 4531 10016 4804 10044
rect 4531 10013 4543 10016
rect 4485 10007 4543 10013
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 4982 10004 4988 10056
rect 5040 10004 5046 10056
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 5810 10044 5816 10056
rect 5767 10016 5816 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5810 10004 5816 10016
rect 5868 10004 5874 10056
rect 6270 10004 6276 10056
rect 6328 10004 6334 10056
rect 6362 10004 6368 10056
rect 6420 10004 6426 10056
rect 10796 10053 10824 10152
rect 11238 10140 11244 10152
rect 11296 10140 11302 10192
rect 11330 10140 11336 10192
rect 11388 10140 11394 10192
rect 11716 10112 11744 10220
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12894 10208 12900 10260
rect 12952 10248 12958 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 12952 10220 14289 10248
rect 12952 10208 12958 10220
rect 14277 10217 14289 10220
rect 14323 10248 14335 10251
rect 14366 10248 14372 10260
rect 14323 10220 14372 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 11072 10084 11744 10112
rect 11072 10053 11100 10084
rect 10781 10047 10839 10053
rect 10781 10013 10793 10047
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 11146 10004 11152 10056
rect 11204 10053 11210 10056
rect 11204 10044 11212 10053
rect 11204 10016 11249 10044
rect 11204 10007 11212 10016
rect 11204 10004 11210 10007
rect 11514 10004 11520 10056
rect 11572 10004 11578 10056
rect 11716 10053 11744 10084
rect 11977 10115 12035 10121
rect 11977 10081 11989 10115
rect 12023 10112 12035 10115
rect 12250 10112 12256 10124
rect 12023 10084 12256 10112
rect 12023 10081 12035 10084
rect 11977 10075 12035 10081
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 16172 10084 16497 10112
rect 16172 10072 16178 10084
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 13354 10004 13360 10056
rect 13412 10004 13418 10056
rect 14734 10044 14740 10056
rect 13556 10016 14740 10044
rect 3082 9948 3556 9976
rect 3620 9948 4200 9976
rect 4249 9979 4307 9985
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 3329 9911 3387 9917
rect 3329 9908 3341 9911
rect 3200 9880 3341 9908
rect 3200 9868 3206 9880
rect 3329 9877 3341 9880
rect 3375 9877 3387 9911
rect 3528 9908 3556 9948
rect 4249 9945 4261 9979
rect 4295 9945 4307 9979
rect 4249 9939 4307 9945
rect 4341 9979 4399 9985
rect 4341 9945 4353 9979
rect 4387 9976 4399 9979
rect 5000 9976 5028 10004
rect 4387 9948 5028 9976
rect 6181 9979 6239 9985
rect 4387 9945 4399 9948
rect 4341 9939 4399 9945
rect 3694 9908 3700 9920
rect 3528 9880 3700 9908
rect 3329 9871 3387 9877
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 4264 9908 4292 9939
rect 4540 9920 4568 9948
rect 6181 9945 6193 9979
rect 6227 9976 6239 9979
rect 6610 9979 6668 9985
rect 6610 9976 6622 9979
rect 6227 9948 6622 9976
rect 6227 9945 6239 9948
rect 6181 9939 6239 9945
rect 6610 9945 6622 9948
rect 6656 9945 6668 9979
rect 6610 9939 6668 9945
rect 10962 9936 10968 9988
rect 11020 9936 11026 9988
rect 11532 9976 11560 10004
rect 12253 9979 12311 9985
rect 11532 9948 11744 9976
rect 4430 9908 4436 9920
rect 4264 9880 4436 9908
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 4522 9868 4528 9920
rect 4580 9868 4586 9920
rect 6270 9868 6276 9920
rect 6328 9908 6334 9920
rect 7742 9908 7748 9920
rect 6328 9880 7748 9908
rect 6328 9868 6334 9880
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 11609 9911 11667 9917
rect 11609 9908 11621 9911
rect 11204 9880 11621 9908
rect 11204 9868 11210 9880
rect 11609 9877 11621 9880
rect 11655 9877 11667 9911
rect 11716 9908 11744 9948
rect 12253 9945 12265 9979
rect 12299 9976 12311 9979
rect 12526 9976 12532 9988
rect 12299 9948 12532 9976
rect 12299 9945 12311 9948
rect 12253 9939 12311 9945
rect 12526 9936 12532 9948
rect 12584 9936 12590 9988
rect 13556 9908 13584 10016
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 14185 9979 14243 9985
rect 14185 9976 14197 9979
rect 13964 9948 14197 9976
rect 13964 9936 13970 9948
rect 14185 9945 14197 9948
rect 14231 9945 14243 9979
rect 14185 9939 14243 9945
rect 15746 9936 15752 9988
rect 15804 9936 15810 9988
rect 11716 9880 13584 9908
rect 11609 9871 11667 9877
rect 13630 9868 13636 9920
rect 13688 9908 13694 9920
rect 13725 9911 13783 9917
rect 13725 9908 13737 9911
rect 13688 9880 13737 9908
rect 13688 9868 13694 9880
rect 13725 9877 13737 9880
rect 13771 9877 13783 9911
rect 13725 9871 13783 9877
rect 14458 9868 14464 9920
rect 14516 9908 14522 9920
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14516 9880 15025 9908
rect 14516 9868 14522 9880
rect 15013 9877 15025 9880
rect 15059 9908 15071 9911
rect 15102 9908 15108 9920
rect 15059 9880 15108 9908
rect 15059 9877 15071 9880
rect 15013 9871 15071 9877
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15838 9868 15844 9920
rect 15896 9908 15902 9920
rect 16776 9908 16804 10007
rect 15896 9880 16804 9908
rect 15896 9868 15902 9880
rect 1104 9818 17112 9840
rect 1104 9766 7214 9818
rect 7266 9766 7278 9818
rect 7330 9766 7342 9818
rect 7394 9766 7406 9818
rect 7458 9766 7470 9818
rect 7522 9766 13214 9818
rect 13266 9766 13278 9818
rect 13330 9766 13342 9818
rect 13394 9766 13406 9818
rect 13458 9766 13470 9818
rect 13522 9766 17112 9818
rect 1104 9744 17112 9766
rect 1854 9664 1860 9716
rect 1912 9704 1918 9716
rect 1949 9707 2007 9713
rect 1949 9704 1961 9707
rect 1912 9676 1961 9704
rect 1912 9664 1918 9676
rect 1949 9673 1961 9676
rect 1995 9673 2007 9707
rect 2774 9704 2780 9716
rect 1949 9667 2007 9673
rect 2700 9676 2780 9704
rect 2700 9636 2728 9676
rect 2774 9664 2780 9676
rect 2832 9664 2838 9716
rect 3050 9664 3056 9716
rect 3108 9664 3114 9716
rect 4522 9664 4528 9716
rect 4580 9664 4586 9716
rect 4614 9664 4620 9716
rect 4672 9664 4678 9716
rect 11238 9664 11244 9716
rect 11296 9664 11302 9716
rect 11330 9664 11336 9716
rect 11388 9664 11394 9716
rect 11885 9707 11943 9713
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 12250 9704 12256 9716
rect 11931 9676 12256 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 12250 9664 12256 9676
rect 12308 9664 12314 9716
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 14182 9704 14188 9716
rect 12584 9676 13032 9704
rect 12584 9664 12590 9676
rect 3068 9636 3096 9664
rect 2056 9608 2728 9636
rect 2792 9608 3096 9636
rect 1854 9528 1860 9580
rect 1912 9528 1918 9580
rect 2056 9577 2084 9608
rect 2792 9577 2820 9608
rect 3694 9596 3700 9648
rect 3752 9596 3758 9648
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9537 2099 9571
rect 2041 9531 2099 9537
rect 2777 9571 2835 9577
rect 2777 9537 2789 9571
rect 2823 9537 2835 9571
rect 4632 9568 4660 9664
rect 8570 9596 8576 9648
rect 8628 9596 8634 9648
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4632 9540 4813 9568
rect 2777 9531 2835 9537
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 10870 9528 10876 9580
rect 10928 9528 10934 9580
rect 11348 9568 11376 9664
rect 13004 9645 13032 9676
rect 13832 9676 14188 9704
rect 12989 9639 13047 9645
rect 12989 9605 13001 9639
rect 13035 9605 13047 9639
rect 13832 9636 13860 9676
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 14826 9664 14832 9716
rect 14884 9704 14890 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14884 9676 14933 9704
rect 14884 9664 14890 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 15838 9704 15844 9716
rect 14921 9667 14979 9673
rect 15396 9676 15844 9704
rect 12989 9599 13047 9605
rect 13188 9608 13860 9636
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11348 9540 11713 9568
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3142 9500 3148 9512
rect 3099 9472 3148 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9469 7711 9503
rect 7653 9463 7711 9469
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 7975 9472 9352 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 7668 9376 7696 9463
rect 4890 9324 4896 9376
rect 4948 9364 4954 9376
rect 4985 9367 5043 9373
rect 4985 9364 4997 9367
rect 4948 9336 4997 9364
rect 4948 9324 4954 9336
rect 4985 9333 4997 9336
rect 5031 9364 5043 9367
rect 6454 9364 6460 9376
rect 5031 9336 6460 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 7650 9324 7656 9376
rect 7708 9324 7714 9376
rect 9324 9364 9352 9472
rect 9490 9460 9496 9512
rect 9548 9460 9554 9512
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9600 9472 9781 9500
rect 9401 9435 9459 9441
rect 9401 9401 9413 9435
rect 9447 9432 9459 9435
rect 9600 9432 9628 9472
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 9447 9404 9628 9432
rect 9447 9401 9459 9404
rect 9401 9395 9459 9401
rect 11146 9364 11152 9376
rect 9324 9336 11152 9364
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 12912 9364 12940 9531
rect 13078 9528 13084 9580
rect 13136 9528 13142 9580
rect 13188 9577 13216 9608
rect 13998 9596 14004 9648
rect 14056 9596 14062 9648
rect 13173 9571 13231 9577
rect 13173 9537 13185 9571
rect 13219 9537 13231 9571
rect 14936 9568 14964 9667
rect 15396 9645 15424 9676
rect 15838 9664 15844 9676
rect 15896 9664 15902 9716
rect 15381 9639 15439 9645
rect 15381 9605 15393 9639
rect 15427 9605 15439 9639
rect 15381 9599 15439 9605
rect 15470 9577 15476 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14936 9540 15025 9568
rect 13173 9531 13231 9537
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9568 15255 9571
rect 15243 9540 15424 9568
rect 15243 9537 15255 9540
rect 15197 9531 15255 9537
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9500 13507 9503
rect 13538 9500 13544 9512
rect 13495 9472 13544 9500
rect 13495 9469 13507 9472
rect 13449 9463 13507 9469
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 15396 9376 15424 9540
rect 15465 9531 15476 9577
rect 15528 9568 15534 9580
rect 15528 9540 15565 9568
rect 15470 9528 15476 9531
rect 15528 9528 15534 9540
rect 14458 9364 14464 9376
rect 12912 9336 14464 9364
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 15010 9324 15016 9376
rect 15068 9324 15074 9376
rect 15378 9324 15384 9376
rect 15436 9324 15442 9376
rect 1104 9274 17112 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 10214 9274
rect 10266 9222 10278 9274
rect 10330 9222 10342 9274
rect 10394 9222 10406 9274
rect 10458 9222 10470 9274
rect 10522 9222 16214 9274
rect 16266 9222 16278 9274
rect 16330 9222 16342 9274
rect 16394 9222 16406 9274
rect 16458 9222 16470 9274
rect 16522 9222 17112 9274
rect 1104 9200 17112 9222
rect 2133 9163 2191 9169
rect 2133 9129 2145 9163
rect 2179 9160 2191 9163
rect 2406 9160 2412 9172
rect 2179 9132 2412 9160
rect 2179 9129 2191 9132
rect 2133 9123 2191 9129
rect 2406 9120 2412 9132
rect 2464 9160 2470 9172
rect 2464 9132 7052 9160
rect 2464 9120 2470 9132
rect 6270 9052 6276 9104
rect 6328 9092 6334 9104
rect 6328 9064 6868 9092
rect 6328 9052 6334 9064
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 9024 4583 9027
rect 4709 9027 4767 9033
rect 4709 9024 4721 9027
rect 4571 8996 4721 9024
rect 4571 8993 4583 8996
rect 4525 8987 4583 8993
rect 4709 8993 4721 8996
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 6512 8996 6776 9024
rect 6512 8984 6518 8996
rect 1854 8956 1860 8968
rect 1596 8928 1860 8956
rect 1596 8832 1624 8928
rect 1854 8916 1860 8928
rect 1912 8956 1918 8968
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1912 8928 2053 8956
rect 1912 8916 1918 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 4632 8888 4660 8919
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 6748 8965 6776 8996
rect 6840 8965 6868 9064
rect 7024 9024 7052 9132
rect 9490 9120 9496 9172
rect 9548 9120 9554 9172
rect 11422 9120 11428 9172
rect 11480 9120 11486 9172
rect 13906 9120 13912 9172
rect 13964 9120 13970 9172
rect 14200 9132 15792 9160
rect 7101 9095 7159 9101
rect 7101 9061 7113 9095
rect 7147 9092 7159 9095
rect 7650 9092 7656 9104
rect 7147 9064 7656 9092
rect 7147 9061 7159 9064
rect 7101 9055 7159 9061
rect 7650 9052 7656 9064
rect 7708 9092 7714 9104
rect 7708 9064 9444 9092
rect 7708 9052 7714 9064
rect 7024 8996 7144 9024
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 6969 8959 7027 8965
rect 6969 8925 6981 8959
rect 7015 8956 7027 8959
rect 7015 8925 7052 8956
rect 6969 8919 7052 8925
rect 4890 8888 4896 8900
rect 4632 8860 4896 8888
rect 4890 8848 4896 8860
rect 4948 8848 4954 8900
rect 4982 8848 4988 8900
rect 5040 8848 5046 8900
rect 1578 8780 1584 8832
rect 1636 8780 1642 8832
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 6564 8820 6592 8919
rect 6512 8792 6592 8820
rect 7024 8820 7052 8919
rect 7116 8888 7144 8996
rect 7742 8984 7748 9036
rect 7800 8984 7806 9036
rect 7653 8959 7711 8965
rect 7653 8925 7665 8959
rect 7699 8956 7711 8959
rect 7760 8956 7788 8984
rect 9416 8965 9444 9064
rect 13357 9027 13415 9033
rect 13357 8993 13369 9027
rect 13403 9024 13415 9027
rect 13630 9024 13636 9036
rect 13403 8996 13636 9024
rect 13403 8993 13415 8996
rect 13357 8987 13415 8993
rect 13630 8984 13636 8996
rect 13688 9024 13694 9036
rect 14200 9024 14228 9132
rect 13688 8996 14228 9024
rect 14645 9027 14703 9033
rect 13688 8984 13694 8996
rect 14645 8993 14657 9027
rect 14691 9024 14703 9027
rect 15010 9024 15016 9036
rect 14691 8996 15016 9024
rect 14691 8993 14703 8996
rect 14645 8987 14703 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 15764 8968 15792 9132
rect 16114 9120 16120 9172
rect 16172 9120 16178 9172
rect 7699 8928 7788 8956
rect 9401 8959 9459 8965
rect 7699 8925 7711 8928
rect 7653 8919 7711 8925
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 10962 8956 10968 8968
rect 9447 8928 10968 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 7116 8860 13032 8888
rect 7558 8820 7564 8832
rect 7024 8792 7564 8820
rect 6512 8780 6518 8792
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 7742 8780 7748 8832
rect 7800 8780 7806 8832
rect 13004 8820 13032 8860
rect 13078 8848 13084 8900
rect 13136 8888 13142 8900
rect 14185 8891 14243 8897
rect 14185 8888 14197 8891
rect 13136 8860 14197 8888
rect 13136 8848 13142 8860
rect 14185 8857 14197 8860
rect 14231 8857 14243 8891
rect 14185 8851 14243 8857
rect 13538 8820 13544 8832
rect 13004 8792 13544 8820
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 14292 8820 14320 8919
rect 14366 8916 14372 8968
rect 14424 8916 14430 8968
rect 15746 8916 15752 8968
rect 15804 8916 15810 8968
rect 15378 8820 15384 8832
rect 14292 8792 15384 8820
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 1104 8730 17112 8752
rect 1104 8678 7214 8730
rect 7266 8678 7278 8730
rect 7330 8678 7342 8730
rect 7394 8678 7406 8730
rect 7458 8678 7470 8730
rect 7522 8678 13214 8730
rect 13266 8678 13278 8730
rect 13330 8678 13342 8730
rect 13394 8678 13406 8730
rect 13458 8678 13470 8730
rect 13522 8678 17112 8730
rect 1104 8656 17112 8678
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5169 8619 5227 8625
rect 5169 8616 5181 8619
rect 5040 8588 5181 8616
rect 5040 8576 5046 8588
rect 5169 8585 5181 8588
rect 5215 8585 5227 8619
rect 5169 8579 5227 8585
rect 7742 8576 7748 8628
rect 7800 8576 7806 8628
rect 13078 8576 13084 8628
rect 13136 8576 13142 8628
rect 13538 8576 13544 8628
rect 13596 8576 13602 8628
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 15470 8616 15476 8628
rect 14424 8588 15476 8616
rect 14424 8576 14430 8588
rect 15470 8576 15476 8588
rect 15528 8616 15534 8628
rect 15528 8588 16528 8616
rect 15528 8576 15534 8588
rect 6086 8548 6092 8560
rect 4922 8520 6092 8548
rect 6086 8508 6092 8520
rect 6144 8508 6150 8560
rect 6365 8551 6423 8557
rect 6365 8517 6377 8551
rect 6411 8548 6423 8551
rect 6454 8548 6460 8560
rect 6411 8520 6460 8548
rect 6411 8517 6423 8520
rect 6365 8511 6423 8517
rect 6454 8508 6460 8520
rect 6512 8508 6518 8560
rect 7024 8520 7604 8548
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3384 8452 3433 8480
rect 3384 8440 3390 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3421 8443 3479 8449
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8480 6055 8483
rect 7024 8480 7052 8520
rect 6043 8452 7052 8480
rect 7101 8483 7159 8489
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8412 3755 8415
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 3743 8384 5917 8412
rect 3743 8381 3755 8384
rect 3697 8375 3755 8381
rect 5905 8381 5917 8384
rect 5951 8381 5963 8415
rect 5905 8375 5963 8381
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7116 8412 7144 8443
rect 7576 8424 7604 8520
rect 7760 8480 7788 8576
rect 8113 8551 8171 8557
rect 8113 8517 8125 8551
rect 8159 8548 8171 8551
rect 8386 8548 8392 8560
rect 8159 8520 8392 8548
rect 8159 8517 8171 8520
rect 8113 8511 8171 8517
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 8570 8508 8576 8560
rect 8628 8508 8634 8560
rect 11333 8551 11391 8557
rect 11333 8517 11345 8551
rect 11379 8548 11391 8551
rect 12989 8551 13047 8557
rect 12989 8548 13001 8551
rect 11379 8520 13001 8548
rect 11379 8517 11391 8520
rect 11333 8511 11391 8517
rect 12989 8517 13001 8520
rect 13035 8517 13047 8551
rect 13096 8548 13124 8576
rect 13096 8520 13492 8548
rect 12989 8511 13047 8517
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7760 8452 7849 8480
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 10928 8452 11161 8480
rect 10928 8440 10934 8452
rect 11149 8449 11161 8452
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11422 8440 11428 8492
rect 11480 8480 11486 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11480 8452 11529 8480
rect 11480 8440 11486 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 13464 8489 13492 8520
rect 13556 8489 13584 8576
rect 16500 8492 16528 8588
rect 11773 8483 11831 8489
rect 11773 8480 11785 8483
rect 11664 8452 11785 8480
rect 11664 8440 11670 8452
rect 11773 8449 11785 8452
rect 11819 8449 11831 8483
rect 11773 8443 11831 8449
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8449 13323 8483
rect 13265 8443 13323 8449
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8449 13507 8483
rect 13449 8443 13507 8449
rect 13541 8483 13599 8489
rect 13541 8449 13553 8483
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 6871 8384 7144 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 7616 8384 9597 8412
rect 7616 8372 7622 8384
rect 9585 8381 9597 8384
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 13280 8412 13308 8443
rect 13722 8440 13728 8492
rect 13780 8440 13786 8492
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 13906 8440 13912 8492
rect 13964 8440 13970 8492
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 16482 8440 16488 8492
rect 16540 8440 16546 8492
rect 13832 8412 13860 8440
rect 13280 8384 13860 8412
rect 5810 8304 5816 8356
rect 5868 8344 5874 8356
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 5868 8316 6653 8344
rect 5868 8304 5874 8316
rect 6641 8313 6653 8316
rect 6687 8313 6699 8347
rect 6641 8307 6699 8313
rect 10965 8347 11023 8353
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 11238 8344 11244 8356
rect 11011 8316 11244 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 11238 8304 11244 8316
rect 11296 8304 11302 8356
rect 12897 8347 12955 8353
rect 12897 8313 12909 8347
rect 12943 8344 12955 8347
rect 13280 8344 13308 8384
rect 15470 8372 15476 8424
rect 15528 8412 15534 8424
rect 16209 8415 16267 8421
rect 16209 8412 16221 8415
rect 15528 8384 16221 8412
rect 15528 8372 15534 8384
rect 16209 8381 16221 8384
rect 16255 8381 16267 8415
rect 16209 8375 16267 8381
rect 12943 8316 13308 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 13354 8304 13360 8356
rect 13412 8304 13418 8356
rect 6914 8236 6920 8288
rect 6972 8236 6978 8288
rect 14550 8236 14556 8288
rect 14608 8236 14614 8288
rect 14734 8236 14740 8288
rect 14792 8236 14798 8288
rect 1104 8186 17112 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 10214 8186
rect 10266 8134 10278 8186
rect 10330 8134 10342 8186
rect 10394 8134 10406 8186
rect 10458 8134 10470 8186
rect 10522 8134 16214 8186
rect 16266 8134 16278 8186
rect 16330 8134 16342 8186
rect 16394 8134 16406 8186
rect 16458 8134 16470 8186
rect 16522 8134 17112 8186
rect 1104 8112 17112 8134
rect 8386 8032 8392 8084
rect 8444 8032 8450 8084
rect 10870 8032 10876 8084
rect 10928 8032 10934 8084
rect 11606 8032 11612 8084
rect 11664 8032 11670 8084
rect 13265 8075 13323 8081
rect 13265 8041 13277 8075
rect 13311 8072 13323 8075
rect 13630 8072 13636 8084
rect 13311 8044 13636 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 14734 8072 14740 8084
rect 13740 8044 14740 8072
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6328 7908 6653 7936
rect 6328 7896 6334 7908
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 6914 7896 6920 7948
rect 6972 7896 6978 7948
rect 3418 7828 3424 7880
rect 3476 7828 3482 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9447 7840 9505 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9493 7837 9505 7840
rect 9539 7868 9551 7871
rect 9582 7868 9588 7880
rect 9539 7840 9588 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 13740 7877 13768 8044
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 14093 7939 14151 7945
rect 14093 7905 14105 7939
rect 14139 7936 14151 7939
rect 14366 7936 14372 7948
rect 14139 7908 14372 7936
rect 14139 7905 14151 7908
rect 14093 7899 14151 7905
rect 14366 7896 14372 7908
rect 14424 7896 14430 7948
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11296 7840 11437 7868
rect 11296 7828 11302 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7868 13507 7871
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13495 7840 13553 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 13814 7828 13820 7880
rect 13872 7828 13878 7880
rect 8570 7800 8576 7812
rect 8142 7772 8576 7800
rect 8220 7744 8248 7772
rect 8570 7760 8576 7772
rect 8628 7760 8634 7812
rect 9766 7809 9772 7812
rect 9760 7763 9772 7809
rect 9766 7760 9772 7763
rect 9824 7760 9830 7812
rect 13173 7803 13231 7809
rect 13173 7769 13185 7803
rect 13219 7800 13231 7803
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 13219 7772 14381 7800
rect 13219 7769 13231 7772
rect 13173 7763 13231 7769
rect 14369 7769 14381 7772
rect 14415 7769 14427 7803
rect 14369 7763 14427 7769
rect 15102 7760 15108 7812
rect 15160 7760 15166 7812
rect 2774 7692 2780 7744
rect 2832 7692 2838 7744
rect 6086 7692 6092 7744
rect 6144 7732 6150 7744
rect 8202 7732 8208 7744
rect 6144 7704 8208 7732
rect 6144 7692 6150 7704
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 15838 7692 15844 7744
rect 15896 7692 15902 7744
rect 1104 7642 17112 7664
rect 1104 7590 7214 7642
rect 7266 7590 7278 7642
rect 7330 7590 7342 7642
rect 7394 7590 7406 7642
rect 7458 7590 7470 7642
rect 7522 7590 13214 7642
rect 13266 7590 13278 7642
rect 13330 7590 13342 7642
rect 13394 7590 13406 7642
rect 13458 7590 13470 7642
rect 13522 7590 17112 7642
rect 1104 7568 17112 7590
rect 2774 7488 2780 7540
rect 2832 7488 2838 7540
rect 4614 7528 4620 7540
rect 4448 7500 4620 7528
rect 2792 7392 2820 7488
rect 4448 7469 4476 7500
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 9766 7488 9772 7540
rect 9824 7488 9830 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11793 7531 11851 7537
rect 11793 7528 11805 7531
rect 11480 7500 11805 7528
rect 11480 7488 11486 7500
rect 11793 7497 11805 7500
rect 11839 7497 11851 7531
rect 11793 7491 11851 7497
rect 13722 7488 13728 7540
rect 13780 7488 13786 7540
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 15470 7528 15476 7540
rect 14783 7500 15476 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 15896 7500 16252 7528
rect 15896 7488 15902 7500
rect 4433 7463 4491 7469
rect 4433 7429 4445 7463
rect 4479 7429 4491 7463
rect 6086 7460 6092 7472
rect 5658 7432 6092 7460
rect 4433 7423 4491 7429
rect 6086 7420 6092 7432
rect 6144 7420 6150 7472
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7460 9367 7463
rect 9355 7432 9996 7460
rect 9355 7429 9367 7432
rect 9309 7423 9367 7429
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2792 7364 2973 7392
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 9490 7352 9496 7404
rect 9548 7352 9554 7404
rect 9674 7352 9680 7404
rect 9732 7352 9738 7404
rect 9968 7401 9996 7432
rect 10962 7420 10968 7472
rect 11020 7460 11026 7472
rect 12710 7460 12716 7472
rect 11020 7432 12716 7460
rect 11020 7420 11026 7432
rect 12710 7420 12716 7432
rect 12768 7420 12774 7472
rect 14185 7463 14243 7469
rect 14185 7429 14197 7463
rect 14231 7460 14243 7463
rect 14550 7460 14556 7472
rect 14231 7432 14556 7460
rect 14231 7429 14243 7432
rect 14185 7423 14243 7429
rect 14550 7420 14556 7432
rect 14608 7420 14614 7472
rect 16224 7469 16252 7500
rect 16209 7463 16267 7469
rect 16209 7429 16221 7463
rect 16255 7429 16267 7463
rect 16209 7423 16267 7429
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 11422 7352 11428 7404
rect 11480 7392 11486 7404
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11480 7364 11989 7392
rect 11480 7352 11486 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 15102 7352 15108 7404
rect 15160 7352 15166 7404
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7392 16543 7395
rect 16574 7392 16580 7404
rect 16531 7364 16580 7392
rect 16531 7361 16543 7364
rect 16485 7355 16543 7361
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 3602 7148 3608 7200
rect 3660 7148 3666 7200
rect 4065 7191 4123 7197
rect 4065 7157 4077 7191
rect 4111 7188 4123 7191
rect 4172 7188 4200 7287
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 15120 7324 15148 7352
rect 15120 7296 16574 7324
rect 16546 7268 16574 7296
rect 16546 7228 16580 7268
rect 16574 7216 16580 7228
rect 16632 7216 16638 7268
rect 4614 7188 4620 7200
rect 4111 7160 4620 7188
rect 4111 7157 4123 7160
rect 4065 7151 4123 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 5905 7191 5963 7197
rect 5905 7157 5917 7191
rect 5951 7188 5963 7191
rect 5994 7188 6000 7200
rect 5951 7160 6000 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 12986 7148 12992 7200
rect 13044 7188 13050 7200
rect 13909 7191 13967 7197
rect 13909 7188 13921 7191
rect 13044 7160 13921 7188
rect 13044 7148 13050 7160
rect 13909 7157 13921 7160
rect 13955 7157 13967 7191
rect 13909 7151 13967 7157
rect 1104 7098 17112 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 10214 7098
rect 10266 7046 10278 7098
rect 10330 7046 10342 7098
rect 10394 7046 10406 7098
rect 10458 7046 10470 7098
rect 10522 7046 16214 7098
rect 16266 7046 16278 7098
rect 16330 7046 16342 7098
rect 16394 7046 16406 7098
rect 16458 7046 16470 7098
rect 16522 7046 17112 7098
rect 1104 7024 17112 7046
rect 5994 6993 6000 6996
rect 5984 6987 6000 6993
rect 5984 6953 5996 6987
rect 5984 6947 6000 6953
rect 5994 6944 6000 6947
rect 6052 6944 6058 6996
rect 9309 6987 9367 6993
rect 9309 6984 9321 6987
rect 8772 6956 9321 6984
rect 7561 6851 7619 6857
rect 7561 6817 7573 6851
rect 7607 6848 7619 6851
rect 7650 6848 7656 6860
rect 7607 6820 7656 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8110 6848 8116 6860
rect 8067 6820 8116 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 8772 6792 8800 6956
rect 9309 6953 9321 6956
rect 9355 6953 9367 6987
rect 9309 6947 9367 6953
rect 9324 6848 9352 6947
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9640 6956 11468 6984
rect 9640 6944 9646 6956
rect 9674 6876 9680 6928
rect 9732 6916 9738 6928
rect 9861 6919 9919 6925
rect 9861 6916 9873 6919
rect 9732 6888 9873 6916
rect 9732 6876 9738 6888
rect 9861 6885 9873 6888
rect 9907 6885 9919 6919
rect 9861 6879 9919 6885
rect 10152 6860 10180 6956
rect 11440 6928 11468 6956
rect 12710 6944 12716 6996
rect 12768 6984 12774 6996
rect 13357 6987 13415 6993
rect 13357 6984 13369 6987
rect 12768 6956 13369 6984
rect 12768 6944 12774 6956
rect 13357 6953 13369 6956
rect 13403 6984 13415 6987
rect 13630 6984 13636 6996
rect 13403 6956 13636 6984
rect 13403 6953 13415 6956
rect 13357 6947 13415 6953
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 16574 6944 16580 6996
rect 16632 6944 16638 6996
rect 11422 6876 11428 6928
rect 11480 6876 11486 6928
rect 12176 6888 12664 6916
rect 8864 6820 9076 6848
rect 9324 6820 9720 6848
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8754 6780 8760 6792
rect 7975 6752 8760 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 5629 6647 5687 6653
rect 5629 6613 5641 6647
rect 5675 6644 5687 6647
rect 5736 6644 5764 6743
rect 8754 6740 8760 6752
rect 8812 6740 8818 6792
rect 8202 6712 8208 6724
rect 7222 6684 8208 6712
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 7006 6644 7012 6656
rect 5675 6616 7012 6644
rect 5675 6613 5687 6616
rect 5629 6607 5687 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 8018 6644 8024 6656
rect 7515 6616 8024 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8864 6644 8892 6820
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 9048 6780 9076 6820
rect 9692 6789 9720 6820
rect 10134 6808 10140 6860
rect 10192 6808 10198 6860
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12176 6857 12204 6888
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 12124 6820 12173 6848
rect 12124 6808 12130 6820
rect 12161 6817 12173 6820
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 12253 6851 12311 6857
rect 12253 6817 12265 6851
rect 12299 6817 12311 6851
rect 12253 6811 12311 6817
rect 9585 6783 9643 6789
rect 9585 6780 9597 6783
rect 9048 6752 9597 6780
rect 8941 6743 8999 6749
rect 9585 6749 9597 6752
rect 9631 6749 9643 6783
rect 9585 6743 9643 6749
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6749 9735 6783
rect 9677 6743 9735 6749
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 12268 6780 12296 6811
rect 12342 6808 12348 6860
rect 12400 6808 12406 6860
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12492 6820 12537 6848
rect 12492 6808 12498 6820
rect 12636 6789 12664 6888
rect 12894 6876 12900 6928
rect 12952 6876 12958 6928
rect 17126 6808 17132 6860
rect 17184 6808 17190 6860
rect 12621 6783 12679 6789
rect 12268 6776 12434 6780
rect 12268 6752 12572 6776
rect 10045 6743 10103 6749
rect 12406 6748 12572 6752
rect 8956 6712 8984 6743
rect 10060 6712 10088 6743
rect 8956 6684 10088 6712
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 8168 6616 9321 6644
rect 8168 6604 8174 6616
rect 9309 6613 9321 6616
rect 9355 6613 9367 6647
rect 9309 6607 9367 6613
rect 9490 6604 9496 6656
rect 9548 6604 9554 6656
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 10060 6644 10088 6684
rect 10410 6672 10416 6724
rect 10468 6672 10474 6724
rect 10962 6672 10968 6724
rect 11020 6672 11026 6724
rect 12544 6712 12572 6748
rect 12621 6749 12633 6783
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6780 12955 6783
rect 13722 6780 13728 6792
rect 12943 6752 13728 6780
rect 12943 6749 12955 6752
rect 12897 6743 12955 6749
rect 12912 6712 12940 6743
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 17144 6780 17172 6808
rect 16807 6752 17172 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 11900 6684 12480 6712
rect 12544 6684 12940 6712
rect 11900 6656 11928 6684
rect 10778 6644 10784 6656
rect 10008 6616 10784 6644
rect 10008 6604 10014 6616
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11882 6604 11888 6656
rect 11940 6604 11946 6656
rect 11974 6604 11980 6656
rect 12032 6604 12038 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 12452 6644 12480 6684
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 13044 6684 13277 6712
rect 13044 6672 13050 6684
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13265 6675 13323 6681
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 12400 6616 12725 6644
rect 12400 6604 12406 6616
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 12713 6607 12771 6613
rect 1104 6554 17112 6576
rect 1104 6502 7214 6554
rect 7266 6502 7278 6554
rect 7330 6502 7342 6554
rect 7394 6502 7406 6554
rect 7458 6502 7470 6554
rect 7522 6502 13214 6554
rect 13266 6502 13278 6554
rect 13330 6502 13342 6554
rect 13394 6502 13406 6554
rect 13458 6502 13470 6554
rect 13522 6502 17112 6554
rect 1104 6480 17112 6502
rect 8754 6400 8760 6452
rect 8812 6400 8818 6452
rect 10045 6443 10103 6449
rect 10045 6409 10057 6443
rect 10091 6440 10103 6443
rect 10134 6440 10140 6452
rect 10091 6412 10140 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 10468 6412 10609 6440
rect 10468 6400 10474 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 11974 6400 11980 6452
rect 12032 6400 12038 6452
rect 12069 6443 12127 6449
rect 12069 6409 12081 6443
rect 12115 6440 12127 6443
rect 12250 6440 12256 6452
rect 12115 6412 12256 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 13817 6443 13875 6449
rect 13817 6409 13829 6443
rect 13863 6409 13875 6443
rect 13817 6403 13875 6409
rect 5166 6372 5172 6384
rect 4724 6344 5172 6372
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 4614 6264 4620 6316
rect 4672 6304 4678 6316
rect 4724 6313 4752 6344
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 7834 6372 7840 6384
rect 7392 6344 7840 6372
rect 4982 6313 4988 6316
rect 4709 6307 4767 6313
rect 4709 6304 4721 6307
rect 4672 6276 4721 6304
rect 4672 6264 4678 6276
rect 4709 6273 4721 6276
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4976 6267 4988 6313
rect 4982 6264 4988 6267
rect 5040 6264 5046 6316
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7392 6313 7420 6344
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 7650 6313 7656 6316
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7064 6276 7297 6304
rect 7064 6264 7070 6276
rect 7285 6273 7297 6276
rect 7331 6304 7343 6307
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7331 6276 7389 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7644 6304 7656 6313
rect 7611 6276 7656 6304
rect 7377 6267 7435 6273
rect 7644 6267 7656 6276
rect 7650 6264 7656 6267
rect 7708 6264 7714 6316
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 11146 6304 11152 6316
rect 10827 6276 11152 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11992 6313 12020 6400
rect 13832 6372 13860 6403
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 15654 6440 15660 6452
rect 13964 6412 15660 6440
rect 13964 6400 13970 6412
rect 14185 6375 14243 6381
rect 14185 6372 14197 6375
rect 13832 6344 14197 6372
rect 14185 6341 14197 6344
rect 14231 6341 14243 6375
rect 14568 6372 14596 6412
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 14568 6344 14674 6372
rect 14185 6335 14243 6341
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6304 12219 6307
rect 12894 6304 12900 6316
rect 12207 6276 12900 6304
rect 12207 6273 12219 6276
rect 12161 6267 12219 6273
rect 12894 6264 12900 6276
rect 12952 6264 12958 6316
rect 13630 6264 13636 6316
rect 13688 6264 13694 6316
rect 2682 6196 2688 6248
rect 2740 6196 2746 6248
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 12250 6236 12256 6248
rect 9548 6208 12256 6236
rect 9548 6196 9554 6208
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6236 13967 6239
rect 13955 6208 13989 6236
rect 13955 6205 13967 6208
rect 13909 6199 13967 6205
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 12986 6168 12992 6180
rect 12216 6140 12992 6168
rect 12216 6128 12222 6140
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 13541 6171 13599 6177
rect 13541 6137 13553 6171
rect 13587 6168 13599 6171
rect 13924 6168 13952 6199
rect 13587 6140 13952 6168
rect 13587 6137 13599 6140
rect 13541 6131 13599 6137
rect 13924 6112 13952 6140
rect 5810 6060 5816 6112
rect 5868 6100 5874 6112
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 5868 6072 6101 6100
rect 5868 6060 5874 6072
rect 6089 6069 6101 6072
rect 6135 6069 6147 6103
rect 6089 6063 6147 6069
rect 13906 6060 13912 6112
rect 13964 6060 13970 6112
rect 14734 6060 14740 6112
rect 14792 6100 14798 6112
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 14792 6072 15669 6100
rect 14792 6060 14798 6072
rect 15657 6069 15669 6072
rect 15703 6069 15715 6103
rect 15657 6063 15715 6069
rect 1104 6010 17112 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 10214 6010
rect 10266 5958 10278 6010
rect 10330 5958 10342 6010
rect 10394 5958 10406 6010
rect 10458 5958 10470 6010
rect 10522 5958 16214 6010
rect 16266 5958 16278 6010
rect 16330 5958 16342 6010
rect 16394 5958 16406 6010
rect 16458 5958 16470 6010
rect 16522 5958 17112 6010
rect 1104 5936 17112 5958
rect 2682 5856 2688 5908
rect 2740 5856 2746 5908
rect 4893 5899 4951 5905
rect 4893 5865 4905 5899
rect 4939 5896 4951 5899
rect 4982 5896 4988 5908
rect 4939 5868 4988 5896
rect 4939 5865 4951 5868
rect 4893 5859 4951 5865
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 10873 5899 10931 5905
rect 10873 5865 10885 5899
rect 10919 5865 10931 5899
rect 10873 5859 10931 5865
rect 2700 5701 2728 5856
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5760 4675 5763
rect 5810 5760 5816 5772
rect 4663 5732 5816 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 9784 5732 10517 5760
rect 9784 5704 9812 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5661 2743 5695
rect 2685 5655 2743 5661
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4890 5692 4896 5704
rect 4571 5664 4896 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 8018 5652 8024 5704
rect 8076 5652 8082 5704
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 9950 5652 9956 5704
rect 10008 5652 10014 5704
rect 10045 5695 10103 5701
rect 10045 5661 10057 5695
rect 10091 5692 10103 5695
rect 10888 5692 10916 5859
rect 11146 5856 11152 5908
rect 11204 5856 11210 5908
rect 13630 5856 13636 5908
rect 13688 5896 13694 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13688 5868 14105 5896
rect 13688 5856 13694 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14093 5859 14151 5865
rect 11793 5763 11851 5769
rect 11793 5729 11805 5763
rect 11839 5760 11851 5763
rect 11882 5760 11888 5772
rect 11839 5732 11888 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 11882 5720 11888 5732
rect 11940 5760 11946 5772
rect 12526 5760 12532 5772
rect 11940 5732 12532 5760
rect 11940 5720 11946 5732
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 14734 5720 14740 5772
rect 14792 5720 14798 5772
rect 10091 5664 10916 5692
rect 11517 5695 11575 5701
rect 10091 5661 10103 5664
rect 10045 5655 10103 5661
rect 11517 5661 11529 5695
rect 11563 5692 11575 5695
rect 12066 5692 12072 5704
rect 11563 5664 12072 5692
rect 11563 5661 11575 5664
rect 11517 5655 11575 5661
rect 3418 5584 3424 5636
rect 3476 5584 3482 5636
rect 8036 5624 8064 5652
rect 10060 5624 10088 5655
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12250 5652 12256 5704
rect 12308 5692 12314 5704
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 12308 5664 12725 5692
rect 12308 5652 12314 5664
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 12860 5664 12909 5692
rect 12860 5652 12866 5664
rect 12897 5661 12909 5664
rect 12943 5692 12955 5695
rect 14461 5695 14519 5701
rect 14461 5692 14473 5695
rect 12943 5664 14473 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 14461 5661 14473 5664
rect 14507 5661 14519 5695
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14461 5655 14519 5661
rect 14752 5664 14933 5692
rect 8036 5596 10088 5624
rect 10413 5627 10471 5633
rect 10413 5593 10425 5627
rect 10459 5593 10471 5627
rect 10413 5587 10471 5593
rect 5166 5516 5172 5568
rect 5224 5516 5230 5568
rect 7745 5559 7803 5565
rect 7745 5525 7757 5559
rect 7791 5556 7803 5559
rect 7834 5556 7840 5568
rect 7791 5528 7840 5556
rect 7791 5525 7803 5528
rect 7745 5519 7803 5525
rect 7834 5516 7840 5528
rect 7892 5556 7898 5568
rect 9582 5556 9588 5568
rect 7892 5528 9588 5556
rect 7892 5516 7898 5528
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 10428 5556 10456 5587
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 10873 5627 10931 5633
rect 10873 5624 10885 5627
rect 10836 5596 10885 5624
rect 10836 5584 10842 5596
rect 10873 5593 10885 5596
rect 10919 5593 10931 5627
rect 12342 5624 12348 5636
rect 10873 5587 10931 5593
rect 10980 5596 12348 5624
rect 10980 5556 11008 5596
rect 12342 5584 12348 5596
rect 12400 5584 12406 5636
rect 13906 5584 13912 5636
rect 13964 5624 13970 5636
rect 14752 5624 14780 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 13964 5596 14780 5624
rect 13964 5584 13970 5596
rect 14752 5568 14780 5596
rect 15194 5584 15200 5636
rect 15252 5584 15258 5636
rect 15654 5584 15660 5636
rect 15712 5584 15718 5636
rect 10428 5528 11008 5556
rect 11054 5516 11060 5568
rect 11112 5516 11118 5568
rect 11606 5516 11612 5568
rect 11664 5516 11670 5568
rect 12805 5559 12863 5565
rect 12805 5525 12817 5559
rect 12851 5556 12863 5559
rect 13814 5556 13820 5568
rect 12851 5528 13820 5556
rect 12851 5525 12863 5528
rect 12805 5519 12863 5525
rect 13814 5516 13820 5528
rect 13872 5556 13878 5568
rect 14553 5559 14611 5565
rect 14553 5556 14565 5559
rect 13872 5528 14565 5556
rect 13872 5516 13878 5528
rect 14553 5525 14565 5528
rect 14599 5525 14611 5559
rect 14553 5519 14611 5525
rect 14734 5516 14740 5568
rect 14792 5516 14798 5568
rect 16666 5516 16672 5568
rect 16724 5516 16730 5568
rect 1104 5466 17112 5488
rect 1104 5414 7214 5466
rect 7266 5414 7278 5466
rect 7330 5414 7342 5466
rect 7394 5414 7406 5466
rect 7458 5414 7470 5466
rect 7522 5414 13214 5466
rect 13266 5414 13278 5466
rect 13330 5414 13342 5466
rect 13394 5414 13406 5466
rect 13458 5414 13470 5466
rect 13522 5414 17112 5466
rect 1104 5392 17112 5414
rect 1578 5312 1584 5364
rect 1636 5312 1642 5364
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 4948 5324 5304 5352
rect 4948 5312 4954 5324
rect 5276 5293 5304 5324
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11793 5355 11851 5361
rect 11793 5352 11805 5355
rect 11112 5324 11805 5352
rect 11112 5312 11118 5324
rect 11793 5321 11805 5324
rect 11839 5352 11851 5355
rect 14277 5355 14335 5361
rect 11839 5324 12434 5352
rect 11839 5321 11851 5324
rect 11793 5315 11851 5321
rect 5261 5287 5319 5293
rect 5261 5253 5273 5287
rect 5307 5284 5319 5287
rect 5537 5287 5595 5293
rect 5537 5284 5549 5287
rect 5307 5256 5549 5284
rect 5307 5253 5319 5256
rect 5261 5247 5319 5253
rect 5537 5253 5549 5256
rect 5583 5284 5595 5287
rect 5626 5284 5632 5296
rect 5583 5256 5632 5284
rect 5583 5253 5595 5256
rect 5537 5247 5595 5253
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 5737 5287 5795 5293
rect 5737 5284 5749 5287
rect 5736 5253 5749 5284
rect 5783 5253 5795 5287
rect 5736 5247 5795 5253
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 992 5188 1409 5216
rect 992 5176 998 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 3780 5219 3838 5225
rect 3780 5185 3792 5219
rect 3826 5216 3838 5219
rect 4062 5216 4068 5228
rect 3826 5188 4068 5216
rect 3826 5185 3838 5188
rect 3780 5179 3838 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5216 5227 5219
rect 5350 5216 5356 5228
rect 5215 5188 5356 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5216 5503 5219
rect 5736 5216 5764 5247
rect 8018 5244 8024 5296
rect 8076 5284 8082 5296
rect 8113 5287 8171 5293
rect 8113 5284 8125 5287
rect 8076 5256 8125 5284
rect 8076 5244 8082 5256
rect 8113 5253 8125 5256
rect 8159 5253 8171 5287
rect 8113 5247 8171 5253
rect 11241 5287 11299 5293
rect 11241 5253 11253 5287
rect 11287 5284 11299 5287
rect 11606 5284 11612 5296
rect 11287 5256 11612 5284
rect 11287 5253 11299 5256
rect 11241 5247 11299 5253
rect 11606 5244 11612 5256
rect 11664 5244 11670 5296
rect 12066 5244 12072 5296
rect 12124 5244 12130 5296
rect 12250 5244 12256 5296
rect 12308 5244 12314 5296
rect 12406 5284 12434 5324
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 15194 5352 15200 5364
rect 14323 5324 15200 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 12621 5287 12679 5293
rect 12621 5284 12633 5287
rect 12406 5256 12633 5284
rect 12621 5253 12633 5256
rect 12667 5284 12679 5287
rect 12802 5284 12808 5296
rect 12667 5256 12808 5284
rect 12667 5253 12679 5256
rect 12621 5247 12679 5253
rect 12802 5244 12808 5256
rect 12860 5244 12866 5296
rect 14553 5287 14611 5293
rect 13648 5256 14228 5284
rect 5491 5188 5764 5216
rect 7009 5219 7067 5225
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 7009 5185 7021 5219
rect 7055 5216 7067 5219
rect 7055 5188 7328 5216
rect 7055 5185 7067 5188
rect 7009 5179 7067 5185
rect 3510 5108 3516 5160
rect 3568 5108 3574 5160
rect 5460 5080 5488 5179
rect 7300 5157 7328 5188
rect 7834 5176 7840 5228
rect 7892 5176 7898 5228
rect 11149 5219 11207 5225
rect 9246 5188 9420 5216
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 7745 5151 7803 5157
rect 7745 5117 7757 5151
rect 7791 5148 7803 5151
rect 8110 5148 8116 5160
rect 7791 5120 8116 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 9392 5148 9420 5188
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11333 5219 11391 5225
rect 11195 5188 11284 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11256 5160 11284 5188
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 11379 5188 11652 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 8260 5120 9420 5148
rect 8260 5108 8266 5120
rect 7469 5083 7527 5089
rect 5460 5052 6776 5080
rect 6748 5024 6776 5052
rect 7469 5049 7481 5083
rect 7515 5080 7527 5083
rect 7558 5080 7564 5092
rect 7515 5052 7564 5080
rect 7515 5049 7527 5052
rect 7469 5043 7527 5049
rect 7558 5040 7564 5052
rect 7616 5040 7622 5092
rect 5258 4972 5264 5024
rect 5316 5012 5322 5024
rect 5445 5015 5503 5021
rect 5445 5012 5457 5015
rect 5316 4984 5457 5012
rect 5316 4972 5322 4984
rect 5445 4981 5457 4984
rect 5491 4981 5503 5015
rect 5445 4975 5503 4981
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5592 4984 5733 5012
rect 5592 4972 5598 4984
rect 5721 4981 5733 4984
rect 5767 5012 5779 5015
rect 5810 5012 5816 5024
rect 5767 4984 5816 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 5905 5015 5963 5021
rect 5905 4981 5917 5015
rect 5951 5012 5963 5015
rect 6362 5012 6368 5024
rect 5951 4984 6368 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6730 4972 6736 5024
rect 6788 4972 6794 5024
rect 7190 4972 7196 5024
rect 7248 4972 7254 5024
rect 9392 5012 9420 5120
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 9766 5148 9772 5160
rect 9631 5120 9772 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 11238 5108 11244 5160
rect 11296 5108 11302 5160
rect 11514 5040 11520 5092
rect 11572 5040 11578 5092
rect 11624 5080 11652 5188
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 11974 5216 11980 5228
rect 11931 5188 11980 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12268 5216 12296 5244
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 12268 5188 12449 5216
rect 12437 5185 12449 5188
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 12820 5148 12848 5244
rect 13648 5225 13676 5256
rect 13814 5225 13820 5228
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 13791 5219 13820 5225
rect 13791 5185 13803 5219
rect 13791 5179 13820 5185
rect 13814 5176 13820 5179
rect 13872 5176 13878 5228
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 13924 5148 13952 5179
rect 13998 5176 14004 5228
rect 14056 5176 14062 5228
rect 14093 5219 14151 5225
rect 14093 5185 14105 5219
rect 14139 5185 14151 5219
rect 14200 5216 14228 5256
rect 14553 5253 14565 5287
rect 14599 5284 14611 5287
rect 14642 5284 14648 5296
rect 14599 5256 14648 5284
rect 14599 5253 14611 5256
rect 14553 5247 14611 5253
rect 14642 5244 14648 5256
rect 14700 5284 14706 5296
rect 16666 5284 16672 5296
rect 14700 5256 14872 5284
rect 14700 5244 14706 5256
rect 14844 5225 14872 5256
rect 16546 5256 16672 5284
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14200 5188 14749 5216
rect 14093 5179 14151 5185
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5185 14887 5219
rect 14829 5179 14887 5185
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5216 15071 5219
rect 16546 5216 16574 5256
rect 16666 5244 16672 5256
rect 16724 5244 16730 5296
rect 15059 5188 16574 5216
rect 15059 5185 15071 5188
rect 15013 5179 15071 5185
rect 12820 5120 13952 5148
rect 14108 5080 14136 5179
rect 14550 5108 14556 5160
rect 14608 5148 14614 5160
rect 14752 5148 14780 5179
rect 15028 5148 15056 5179
rect 14608 5120 15056 5148
rect 14608 5108 14614 5120
rect 14369 5083 14427 5089
rect 14369 5080 14381 5083
rect 11624 5052 12296 5080
rect 12158 5012 12164 5024
rect 9392 4984 12164 5012
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 12268 5021 12296 5052
rect 13280 5052 14381 5080
rect 13280 5024 13308 5052
rect 14369 5049 14381 5052
rect 14415 5049 14427 5083
rect 14369 5043 14427 5049
rect 12253 5015 12311 5021
rect 12253 4981 12265 5015
rect 12299 5012 12311 5015
rect 12986 5012 12992 5024
rect 12299 4984 12992 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 13262 4972 13268 5024
rect 13320 4972 13326 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14458 5012 14464 5024
rect 14056 4984 14464 5012
rect 14056 4972 14062 4984
rect 14458 4972 14464 4984
rect 14516 5012 14522 5024
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 14516 4984 14933 5012
rect 14516 4972 14522 4984
rect 14921 4981 14933 4984
rect 14967 4981 14979 5015
rect 14921 4975 14979 4981
rect 1104 4922 17112 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 10214 4922
rect 10266 4870 10278 4922
rect 10330 4870 10342 4922
rect 10394 4870 10406 4922
rect 10458 4870 10470 4922
rect 10522 4870 16214 4922
rect 16266 4870 16278 4922
rect 16330 4870 16342 4922
rect 16394 4870 16406 4922
rect 16458 4870 16470 4922
rect 16522 4870 17112 4922
rect 1104 4848 17112 4870
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 4120 4780 4169 4808
rect 4120 4768 4126 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 5626 4808 5632 4820
rect 4157 4771 4215 4777
rect 4264 4780 5632 4808
rect 4264 4613 4292 4780
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 8202 4808 8208 4820
rect 7064 4780 8208 4808
rect 7064 4768 7070 4780
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 9217 4811 9275 4817
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9582 4808 9588 4820
rect 9263 4780 9588 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 5166 4672 5172 4684
rect 5031 4644 5172 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5166 4632 5172 4644
rect 5224 4672 5230 4684
rect 9324 4681 9352 4780
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 11238 4768 11244 4820
rect 11296 4768 11302 4820
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 12713 4811 12771 4817
rect 12713 4808 12725 4811
rect 11572 4780 12725 4808
rect 11572 4768 11578 4780
rect 12713 4777 12725 4780
rect 12759 4777 12771 4811
rect 12713 4771 12771 4777
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13446 4808 13452 4820
rect 13403 4780 13452 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 11149 4743 11207 4749
rect 11149 4709 11161 4743
rect 11195 4709 11207 4743
rect 11149 4703 11207 4709
rect 11256 4740 11284 4768
rect 11885 4743 11943 4749
rect 11885 4740 11897 4743
rect 11256 4712 11897 4740
rect 9309 4675 9367 4681
rect 5224 4644 5396 4672
rect 5224 4632 5230 4644
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5092 4468 5120 4567
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 5368 4613 5396 4644
rect 9309 4641 9321 4675
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 11164 4672 11192 4703
rect 9631 4644 11192 4672
rect 11256 4672 11284 4712
rect 11885 4709 11897 4712
rect 11931 4709 11943 4743
rect 11885 4703 11943 4709
rect 11256 4644 11468 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 7098 4604 7104 4616
rect 5399 4576 7104 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 7098 4564 7104 4576
rect 7156 4604 7162 4616
rect 7834 4604 7840 4616
rect 7156 4576 7840 4604
rect 7156 4564 7162 4576
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 10962 4604 10968 4616
rect 10718 4576 10968 4604
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11330 4564 11336 4616
rect 11388 4564 11394 4616
rect 11440 4613 11468 4644
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 11664 4644 11805 4672
rect 11664 4632 11670 4644
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 11793 4635 11851 4641
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 12032 4644 12081 4672
rect 12032 4632 12038 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12621 4675 12679 4681
rect 12621 4672 12633 4675
rect 12069 4635 12127 4641
rect 12176 4644 12633 4672
rect 12176 4613 12204 4644
rect 12621 4641 12633 4644
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4573 11483 4607
rect 11425 4567 11483 4573
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 5169 4539 5227 4545
rect 5169 4505 5181 4539
rect 5215 4536 5227 4539
rect 5598 4539 5656 4545
rect 5598 4536 5610 4539
rect 5215 4508 5610 4536
rect 5215 4505 5227 4508
rect 5169 4499 5227 4505
rect 5598 4505 5610 4508
rect 5644 4505 5656 4539
rect 5598 4499 5656 4505
rect 6362 4496 6368 4548
rect 6420 4496 6426 4548
rect 7190 4496 7196 4548
rect 7248 4536 7254 4548
rect 7346 4539 7404 4545
rect 7346 4536 7358 4539
rect 7248 4508 7358 4536
rect 7248 4496 7254 4508
rect 7346 4505 7358 4508
rect 7392 4505 7404 4539
rect 11698 4536 11704 4548
rect 7346 4499 7404 4505
rect 11072 4508 11704 4536
rect 6380 4468 6408 4496
rect 5092 4440 6408 4468
rect 6730 4428 6736 4480
rect 6788 4428 6794 4480
rect 8478 4428 8484 4480
rect 8536 4428 8542 4480
rect 11072 4477 11100 4508
rect 11698 4496 11704 4508
rect 11756 4536 11762 4548
rect 12176 4536 12204 4567
rect 11756 4508 12204 4536
rect 12268 4536 12296 4567
rect 12342 4564 12348 4616
rect 12400 4564 12406 4616
rect 12526 4564 12532 4616
rect 12584 4564 12590 4616
rect 12728 4536 12756 4771
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 13538 4768 13544 4820
rect 13596 4768 13602 4820
rect 14277 4811 14335 4817
rect 14277 4777 14289 4811
rect 14323 4808 14335 4811
rect 14550 4808 14556 4820
rect 14323 4780 14556 4808
rect 14323 4777 14335 4780
rect 14277 4771 14335 4777
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 13262 4632 13268 4684
rect 13320 4632 13326 4684
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4604 12863 4607
rect 12894 4604 12900 4616
rect 12851 4576 12900 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4604 13415 4607
rect 13403 4576 14228 4604
rect 13403 4573 13415 4576
rect 13357 4567 13415 4573
rect 13081 4539 13139 4545
rect 13081 4536 13093 4539
rect 12268 4508 12756 4536
rect 13004 4508 13093 4536
rect 11756 4496 11762 4508
rect 13004 4477 13032 4508
rect 13081 4505 13093 4508
rect 13127 4505 13139 4539
rect 13081 4499 13139 4505
rect 11057 4471 11115 4477
rect 11057 4437 11069 4471
rect 11103 4437 11115 4471
rect 11057 4431 11115 4437
rect 12989 4471 13047 4477
rect 12989 4437 13001 4471
rect 13035 4437 13047 4471
rect 12989 4431 13047 4437
rect 13906 4428 13912 4480
rect 13964 4468 13970 4480
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 13964 4440 14105 4468
rect 13964 4428 13970 4440
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14200 4468 14228 4576
rect 14461 4539 14519 4545
rect 14461 4505 14473 4539
rect 14507 4536 14519 4539
rect 14642 4536 14648 4548
rect 14507 4508 14648 4536
rect 14507 4505 14519 4508
rect 14461 4499 14519 4505
rect 14642 4496 14648 4508
rect 14700 4496 14706 4548
rect 14274 4477 14280 4480
rect 14261 4471 14280 4477
rect 14261 4468 14273 4471
rect 14200 4440 14273 4468
rect 14093 4431 14151 4437
rect 14261 4437 14273 4440
rect 14261 4431 14280 4437
rect 14274 4428 14280 4431
rect 14332 4428 14338 4480
rect 14734 4428 14740 4480
rect 14792 4428 14798 4480
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15562 4468 15568 4480
rect 15252 4440 15568 4468
rect 15252 4428 15258 4440
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 1104 4378 17112 4400
rect 1104 4326 7214 4378
rect 7266 4326 7278 4378
rect 7330 4326 7342 4378
rect 7394 4326 7406 4378
rect 7458 4326 7470 4378
rect 7522 4326 13214 4378
rect 13266 4326 13278 4378
rect 13330 4326 13342 4378
rect 13394 4326 13406 4378
rect 13458 4326 13470 4378
rect 13522 4326 17112 4378
rect 1104 4304 17112 4326
rect 5810 4224 5816 4276
rect 5868 4224 5874 4276
rect 5997 4267 6055 4273
rect 5997 4233 6009 4267
rect 6043 4264 6055 4267
rect 6730 4264 6736 4276
rect 6043 4236 6736 4264
rect 6043 4233 6055 4236
rect 5997 4227 6055 4233
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7098 4264 7104 4276
rect 7055 4236 7104 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7469 4267 7527 4273
rect 7469 4233 7481 4267
rect 7515 4264 7527 4267
rect 7558 4264 7564 4276
rect 7515 4236 7564 4264
rect 7515 4233 7527 4236
rect 7469 4227 7527 4233
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 8297 4267 8355 4273
rect 8297 4264 8309 4267
rect 7852 4236 8309 4264
rect 3237 4199 3295 4205
rect 3237 4196 3249 4199
rect 2746 4168 3249 4196
rect 14 4088 20 4140
rect 72 4128 78 4140
rect 2746 4128 2774 4168
rect 3237 4165 3249 4168
rect 3283 4196 3295 4199
rect 3418 4196 3424 4208
rect 3283 4168 3424 4196
rect 3283 4165 3295 4168
rect 3237 4159 3295 4165
rect 3418 4156 3424 4168
rect 3476 4156 3482 4208
rect 3510 4156 3516 4208
rect 3568 4196 3574 4208
rect 4065 4199 4123 4205
rect 4065 4196 4077 4199
rect 3568 4168 4077 4196
rect 3568 4156 3574 4168
rect 4065 4165 4077 4168
rect 4111 4196 4123 4199
rect 5166 4196 5172 4208
rect 4111 4168 5172 4196
rect 4111 4165 4123 4168
rect 4065 4159 4123 4165
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 5626 4156 5632 4208
rect 5684 4156 5690 4208
rect 5905 4199 5963 4205
rect 5905 4165 5917 4199
rect 5951 4196 5963 4199
rect 6270 4196 6276 4208
rect 5951 4168 6276 4196
rect 5951 4165 5963 4168
rect 5905 4159 5963 4165
rect 6270 4156 6276 4168
rect 6328 4196 6334 4208
rect 6328 4168 6592 4196
rect 6328 4156 6334 4168
rect 72 4100 2774 4128
rect 72 4088 78 4100
rect 6362 4088 6368 4140
rect 6420 4088 6426 4140
rect 6564 4137 6592 4168
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 7852 4128 7880 4236
rect 8297 4233 8309 4236
rect 8343 4233 8355 4267
rect 8297 4227 8355 4233
rect 8389 4267 8447 4273
rect 8389 4233 8401 4267
rect 8435 4264 8447 4267
rect 8478 4264 8484 4276
rect 8435 4236 8484 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 8110 4156 8116 4208
rect 8168 4156 8174 4208
rect 8404 4196 8432 4227
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 11057 4267 11115 4273
rect 11057 4233 11069 4267
rect 11103 4264 11115 4267
rect 11330 4264 11336 4276
rect 11103 4236 11336 4264
rect 11103 4233 11115 4236
rect 11057 4227 11115 4233
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 13630 4264 13636 4276
rect 12636 4236 13636 4264
rect 8220 4168 8432 4196
rect 6549 4091 6607 4097
rect 7668 4100 7880 4128
rect 7929 4131 7987 4137
rect 7668 4069 7696 4100
rect 7929 4097 7941 4131
rect 7975 4128 7987 4131
rect 8220 4128 8248 4168
rect 11514 4156 11520 4208
rect 11572 4156 11578 4208
rect 7975 4100 8248 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 8478 4088 8484 4140
rect 8536 4088 8542 4140
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4128 11115 4131
rect 11146 4128 11152 4140
rect 11103 4100 11152 4128
rect 11103 4097 11115 4100
rect 11057 4091 11115 4097
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 6472 4032 7665 4060
rect 6472 4004 6500 4032
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 8202 4060 8208 4072
rect 7883 4032 8208 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 6181 3995 6239 4001
rect 6181 3961 6193 3995
rect 6227 3992 6239 3995
rect 6454 3992 6460 4004
rect 6227 3964 6460 3992
rect 6227 3961 6239 3964
rect 6181 3955 6239 3961
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 7760 3992 7788 4023
rect 8202 4020 8208 4032
rect 8260 4060 8266 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 8260 4032 8677 4060
rect 8260 4020 8266 4032
rect 8665 4029 8677 4032
rect 8711 4029 8723 4063
rect 10888 4060 10916 4091
rect 11146 4088 11152 4100
rect 11204 4128 11210 4140
rect 11532 4128 11560 4156
rect 11204 4100 11560 4128
rect 11204 4088 11210 4100
rect 11606 4088 11612 4140
rect 11664 4128 11670 4140
rect 12342 4128 12348 4140
rect 11664 4100 12348 4128
rect 11664 4088 11670 4100
rect 12342 4088 12348 4100
rect 12400 4128 12406 4140
rect 12636 4137 12664 4236
rect 13630 4224 13636 4236
rect 13688 4264 13694 4276
rect 13688 4236 13768 4264
rect 13688 4224 13694 4236
rect 12710 4156 12716 4208
rect 12768 4196 12774 4208
rect 13538 4196 13544 4208
rect 12768 4168 13544 4196
rect 12768 4156 12774 4168
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 13740 4205 13768 4236
rect 13725 4199 13783 4205
rect 13725 4165 13737 4199
rect 13771 4165 13783 4199
rect 13725 4159 13783 4165
rect 13906 4156 13912 4208
rect 13964 4156 13970 4208
rect 14093 4199 14151 4205
rect 14093 4165 14105 4199
rect 14139 4196 14151 4199
rect 14274 4196 14280 4208
rect 14139 4168 14280 4196
rect 14139 4165 14151 4168
rect 14093 4159 14151 4165
rect 14274 4156 14280 4168
rect 14332 4196 14338 4208
rect 14332 4168 14596 4196
rect 14332 4156 14338 4168
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12400 4100 12633 4128
rect 12400 4088 12406 4100
rect 12621 4097 12633 4100
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4097 12863 4131
rect 12805 4091 12863 4097
rect 11422 4060 11428 4072
rect 10888 4032 11428 4060
rect 8665 4023 8723 4029
rect 11422 4020 11428 4032
rect 11480 4060 11486 4072
rect 11974 4060 11980 4072
rect 11480 4032 11980 4060
rect 11480 4020 11486 4032
rect 11974 4020 11980 4032
rect 12032 4060 12038 4072
rect 12820 4060 12848 4091
rect 12986 4088 12992 4140
rect 13044 4128 13050 4140
rect 13265 4131 13323 4137
rect 13265 4128 13277 4131
rect 13044 4100 13277 4128
rect 13044 4088 13050 4100
rect 13265 4097 13277 4100
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4128 13507 4131
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 13495 4100 14381 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13357 4063 13415 4069
rect 12032 4032 13032 4060
rect 12032 4020 12038 4032
rect 8478 3992 8484 4004
rect 7760 3964 8484 3992
rect 8478 3952 8484 3964
rect 8536 3952 8542 4004
rect 13004 3936 13032 4032
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 13998 4060 14004 4072
rect 13403 4032 14004 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 13541 3995 13599 4001
rect 13541 3961 13553 3995
rect 13587 3992 13599 3995
rect 14108 3992 14136 4100
rect 14369 4097 14381 4100
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14458 4088 14464 4140
rect 14516 4088 14522 4140
rect 13587 3964 14136 3992
rect 13587 3961 13599 3964
rect 13541 3955 13599 3961
rect 6362 3884 6368 3936
rect 6420 3884 6426 3936
rect 12802 3884 12808 3936
rect 12860 3884 12866 3936
rect 12986 3884 12992 3936
rect 13044 3884 13050 3936
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 13906 3924 13912 3936
rect 13228 3896 13912 3924
rect 13228 3884 13234 3896
rect 13906 3884 13912 3896
rect 13964 3884 13970 3936
rect 14568 3924 14596 4168
rect 15562 4156 15568 4208
rect 15620 4156 15626 4208
rect 14734 4088 14740 4140
rect 14792 4088 14798 4140
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 14660 4032 15025 4060
rect 14660 4001 14688 4032
rect 15013 4029 15025 4032
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 14645 3995 14703 4001
rect 14645 3961 14657 3995
rect 14691 3961 14703 3995
rect 14645 3955 14703 3961
rect 16485 3927 16543 3933
rect 16485 3924 16497 3927
rect 14568 3896 16497 3924
rect 16485 3893 16497 3896
rect 16531 3893 16543 3927
rect 16485 3887 16543 3893
rect 1104 3834 17112 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 10214 3834
rect 10266 3782 10278 3834
rect 10330 3782 10342 3834
rect 10394 3782 10406 3834
rect 10458 3782 10470 3834
rect 10522 3782 16214 3834
rect 16266 3782 16278 3834
rect 16330 3782 16342 3834
rect 16394 3782 16406 3834
rect 16458 3782 16470 3834
rect 16522 3782 17112 3834
rect 1104 3760 17112 3782
rect 4801 3723 4859 3729
rect 4801 3689 4813 3723
rect 4847 3720 4859 3723
rect 5166 3720 5172 3732
rect 4847 3692 5172 3720
rect 4847 3689 4859 3692
rect 4801 3683 4859 3689
rect 4908 3593 4936 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 6270 3680 6276 3732
rect 6328 3680 6334 3732
rect 6362 3680 6368 3732
rect 6420 3680 6426 3732
rect 6454 3680 6460 3732
rect 6512 3680 6518 3732
rect 12802 3720 12808 3732
rect 12452 3692 12808 3720
rect 4893 3587 4951 3593
rect 4893 3553 4905 3587
rect 4939 3553 4951 3587
rect 4893 3547 4951 3553
rect 6380 3525 6408 3680
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6472 3516 6500 3680
rect 7668 3624 8708 3652
rect 7668 3525 7696 3624
rect 8478 3584 8484 3596
rect 7852 3556 8484 3584
rect 7852 3525 7880 3556
rect 8478 3544 8484 3556
rect 8536 3584 8542 3596
rect 8536 3556 8616 3584
rect 8536 3544 8542 3556
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6472 3488 6561 3516
rect 6365 3479 6423 3485
rect 6549 3485 6561 3488
rect 6595 3516 6607 3519
rect 7653 3519 7711 3525
rect 7653 3516 7665 3519
rect 6595 3488 7665 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 7653 3485 7665 3488
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3516 8079 3519
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8067 3488 8309 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8588 3525 8616 3556
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8680 3516 8708 3624
rect 11072 3556 12388 3584
rect 11072 3525 11100 3556
rect 8757 3519 8815 3525
rect 8757 3516 8769 3519
rect 8680 3488 8769 3516
rect 8573 3479 8631 3485
rect 8757 3485 8769 3488
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 11146 3476 11152 3528
rect 11204 3476 11210 3528
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 11514 3476 11520 3528
rect 11572 3476 11578 3528
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 5160 3451 5218 3457
rect 5160 3417 5172 3451
rect 5206 3448 5218 3451
rect 6457 3451 6515 3457
rect 6457 3448 6469 3451
rect 5206 3420 6469 3448
rect 5206 3417 5218 3420
rect 5160 3411 5218 3417
rect 6457 3417 6469 3420
rect 6503 3417 6515 3451
rect 8404 3448 8432 3476
rect 8665 3451 8723 3457
rect 8665 3448 8677 3451
rect 8404 3420 8677 3448
rect 6457 3411 6515 3417
rect 8665 3417 8677 3420
rect 8711 3417 8723 3451
rect 8665 3411 8723 3417
rect 8110 3340 8116 3392
rect 8168 3340 8174 3392
rect 10134 3340 10140 3392
rect 10192 3380 10198 3392
rect 10873 3383 10931 3389
rect 10873 3380 10885 3383
rect 10192 3352 10885 3380
rect 10192 3340 10198 3352
rect 10873 3349 10885 3352
rect 10919 3349 10931 3383
rect 11164 3380 11192 3476
rect 11241 3451 11299 3457
rect 11241 3417 11253 3451
rect 11287 3448 11299 3451
rect 11609 3451 11667 3457
rect 11609 3448 11621 3451
rect 11287 3420 11621 3448
rect 11287 3417 11299 3420
rect 11241 3411 11299 3417
rect 11609 3417 11621 3420
rect 11655 3417 11667 3451
rect 11609 3411 11667 3417
rect 11716 3380 11744 3479
rect 11164 3352 11744 3380
rect 10873 3343 10931 3349
rect 12066 3340 12072 3392
rect 12124 3380 12130 3392
rect 12253 3383 12311 3389
rect 12253 3380 12265 3383
rect 12124 3352 12265 3380
rect 12124 3340 12130 3352
rect 12253 3349 12265 3352
rect 12299 3349 12311 3383
rect 12360 3380 12388 3556
rect 12452 3525 12480 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 13173 3723 13231 3729
rect 13173 3720 13185 3723
rect 12952 3692 13185 3720
rect 12952 3680 12958 3692
rect 13173 3689 13185 3692
rect 13219 3689 13231 3723
rect 13173 3683 13231 3689
rect 13998 3680 14004 3732
rect 14056 3680 14062 3732
rect 13078 3652 13084 3664
rect 12544 3624 13084 3652
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 12544 3457 12572 3624
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 12802 3544 12808 3596
rect 12860 3584 12866 3596
rect 14016 3584 14044 3680
rect 12860 3556 13400 3584
rect 14016 3556 14504 3584
rect 12860 3544 12866 3556
rect 12894 3476 12900 3528
rect 12952 3476 12958 3528
rect 13372 3518 13400 3556
rect 13449 3519 13507 3525
rect 13449 3518 13461 3519
rect 13004 3488 13308 3516
rect 13372 3490 13461 3518
rect 12529 3451 12587 3457
rect 12529 3417 12541 3451
rect 12575 3417 12587 3451
rect 12529 3411 12587 3417
rect 12618 3408 12624 3460
rect 12676 3408 12682 3460
rect 12739 3451 12797 3457
rect 12739 3448 12751 3451
rect 12728 3417 12751 3448
rect 12785 3448 12797 3451
rect 13004 3448 13032 3488
rect 12785 3420 13032 3448
rect 12785 3417 12797 3420
rect 12728 3411 12797 3417
rect 12728 3380 12756 3411
rect 12360 3352 12756 3380
rect 12253 3343 12311 3349
rect 12986 3340 12992 3392
rect 13044 3340 13050 3392
rect 13170 3389 13176 3392
rect 13157 3383 13176 3389
rect 13157 3349 13169 3383
rect 13157 3343 13176 3349
rect 13170 3340 13176 3343
rect 13228 3340 13234 3392
rect 13280 3380 13308 3488
rect 13449 3485 13461 3490
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3510 13691 3519
rect 13722 3510 13728 3528
rect 13679 3485 13728 3510
rect 13633 3482 13728 3485
rect 13633 3479 13691 3482
rect 13722 3476 13728 3482
rect 13780 3476 13786 3528
rect 13906 3476 13912 3528
rect 13964 3516 13970 3528
rect 14476 3525 14504 3556
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13964 3488 14105 3516
rect 13964 3476 13970 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 14093 3479 14151 3485
rect 14200 3488 14381 3516
rect 13357 3451 13415 3457
rect 13357 3417 13369 3451
rect 13403 3448 13415 3451
rect 13538 3448 13544 3460
rect 13403 3420 13544 3448
rect 13403 3417 13415 3420
rect 13357 3411 13415 3417
rect 13538 3408 13544 3420
rect 13596 3448 13602 3460
rect 14200 3448 14228 3488
rect 14369 3485 14381 3488
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 13596 3420 14228 3448
rect 13596 3408 13602 3420
rect 14274 3408 14280 3460
rect 14332 3408 14338 3460
rect 13817 3383 13875 3389
rect 13817 3380 13829 3383
rect 13280 3352 13829 3380
rect 13817 3349 13829 3352
rect 13863 3349 13875 3383
rect 13817 3343 13875 3349
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 15286 3380 15292 3392
rect 14691 3352 15292 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 1104 3290 17112 3312
rect 1104 3238 7214 3290
rect 7266 3238 7278 3290
rect 7330 3238 7342 3290
rect 7394 3238 7406 3290
rect 7458 3238 7470 3290
rect 7522 3238 13214 3290
rect 13266 3238 13278 3290
rect 13330 3238 13342 3290
rect 13394 3238 13406 3290
rect 13458 3238 13470 3290
rect 13522 3238 17112 3290
rect 1104 3216 17112 3238
rect 7098 3136 7104 3188
rect 7156 3136 7162 3188
rect 8021 3179 8079 3185
rect 8021 3145 8033 3179
rect 8067 3176 8079 3179
rect 8478 3176 8484 3188
rect 8067 3148 8484 3176
rect 8067 3145 8079 3148
rect 8021 3139 8079 3145
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 11698 3176 11704 3188
rect 9640 3148 11704 3176
rect 9640 3136 9646 3148
rect 6181 3111 6239 3117
rect 6181 3077 6193 3111
rect 6227 3108 6239 3111
rect 7116 3108 7144 3136
rect 6227 3080 7144 3108
rect 6227 3077 6239 3080
rect 6181 3071 6239 3077
rect 6656 3049 6684 3080
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 6908 3043 6966 3049
rect 6908 3009 6920 3043
rect 6954 3040 6966 3043
rect 7190 3040 7196 3052
rect 6954 3012 7196 3040
rect 6954 3009 6966 3012
rect 6908 3003 6966 3009
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 9600 3049 9628 3136
rect 9861 3111 9919 3117
rect 9861 3077 9873 3111
rect 9907 3108 9919 3111
rect 10134 3108 10140 3120
rect 9907 3080 10140 3108
rect 9907 3077 9919 3080
rect 9861 3071 9919 3077
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 9226 3043 9284 3049
rect 9226 3040 9238 3043
rect 8536 3012 9238 3040
rect 8536 3000 8542 3012
rect 9226 3009 9238 3012
rect 9272 3009 9284 3043
rect 9226 3003 9284 3009
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3040 9551 3043
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 9539 3012 9597 3040
rect 9539 3009 9551 3012
rect 9493 3003 9551 3009
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 10962 3000 10968 3052
rect 11020 3000 11026 3052
rect 11532 3049 11560 3148
rect 11698 3136 11704 3148
rect 11756 3176 11762 3188
rect 13633 3179 13691 3185
rect 13633 3176 13645 3179
rect 11756 3148 13645 3176
rect 11756 3136 11762 3148
rect 13633 3145 13645 3148
rect 13679 3176 13691 3179
rect 14734 3176 14740 3188
rect 13679 3148 14740 3176
rect 13679 3145 13691 3148
rect 13633 3139 13691 3145
rect 14734 3136 14740 3148
rect 14792 3176 14798 3188
rect 14792 3148 15884 3176
rect 14792 3136 14798 3148
rect 11793 3111 11851 3117
rect 11793 3077 11805 3111
rect 11839 3108 11851 3111
rect 12066 3108 12072 3120
rect 11839 3080 12072 3108
rect 11839 3077 11851 3080
rect 11793 3071 11851 3077
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 13817 3111 13875 3117
rect 13817 3077 13829 3111
rect 13863 3108 13875 3111
rect 14274 3108 14280 3120
rect 13863 3080 14280 3108
rect 13863 3077 13875 3080
rect 13817 3071 13875 3077
rect 14274 3068 14280 3080
rect 14332 3068 14338 3120
rect 15102 3068 15108 3120
rect 15160 3068 15166 3120
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 15565 3111 15623 3117
rect 15565 3108 15577 3111
rect 15344 3080 15577 3108
rect 15344 3068 15350 3080
rect 15565 3077 15577 3080
rect 15611 3077 15623 3111
rect 15565 3071 15623 3077
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 10980 2972 11008 3000
rect 12912 2972 12940 3026
rect 13538 3000 13544 3052
rect 13596 3000 13602 3052
rect 13630 3000 13636 3052
rect 13688 3040 13694 3052
rect 15856 3049 15884 3148
rect 13725 3043 13783 3049
rect 13725 3040 13737 3043
rect 13688 3012 13737 3040
rect 13688 3000 13694 3012
rect 13725 3009 13737 3012
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 10980 2944 12940 2972
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13265 2975 13323 2981
rect 13265 2972 13277 2975
rect 13044 2944 13277 2972
rect 13044 2932 13050 2944
rect 13265 2941 13277 2944
rect 13311 2941 13323 2975
rect 13556 2972 13584 3000
rect 13924 2972 13952 3003
rect 14093 2975 14151 2981
rect 14093 2972 14105 2975
rect 13556 2944 14105 2972
rect 13265 2935 13323 2941
rect 14093 2941 14105 2944
rect 14139 2941 14151 2975
rect 14093 2935 14151 2941
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 11333 2907 11391 2913
rect 11333 2904 11345 2907
rect 11204 2876 11345 2904
rect 11204 2864 11210 2876
rect 11333 2873 11345 2876
rect 11379 2873 11391 2907
rect 11333 2867 11391 2873
rect 8113 2839 8171 2845
rect 8113 2805 8125 2839
rect 8159 2836 8171 2839
rect 8202 2836 8208 2848
rect 8159 2808 8208 2836
rect 8159 2805 8171 2808
rect 8113 2799 8171 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 1104 2746 17112 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 10214 2746
rect 10266 2694 10278 2746
rect 10330 2694 10342 2746
rect 10394 2694 10406 2746
rect 10458 2694 10470 2746
rect 10522 2694 16214 2746
rect 16266 2694 16278 2746
rect 16330 2694 16342 2746
rect 16394 2694 16406 2746
rect 16458 2694 16470 2746
rect 16522 2694 17112 2746
rect 1104 2672 17112 2694
rect 7190 2592 7196 2644
rect 7248 2592 7254 2644
rect 7837 2635 7895 2641
rect 7837 2601 7849 2635
rect 7883 2632 7895 2635
rect 9490 2632 9496 2644
rect 7883 2604 9496 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10594 2632 10600 2644
rect 9999 2604 10600 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 11698 2592 11704 2644
rect 11756 2592 11762 2644
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 16301 2635 16359 2641
rect 16301 2632 16313 2635
rect 15436 2604 16313 2632
rect 15436 2592 15442 2604
rect 16301 2601 16313 2604
rect 16347 2601 16359 2635
rect 16301 2595 16359 2601
rect 8110 2564 8116 2576
rect 7392 2536 8116 2564
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2428 4859 2431
rect 7006 2428 7012 2440
rect 4847 2400 7012 2428
rect 4847 2397 4859 2400
rect 4801 2391 4859 2397
rect 7006 2388 7012 2400
rect 7064 2388 7070 2440
rect 7392 2437 7420 2536
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 8478 2524 8484 2576
rect 8536 2524 8542 2576
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 8386 2496 8392 2508
rect 8251 2468 8392 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 8159 2400 8248 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 8220 2372 8248 2400
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2428 16543 2431
rect 17034 2428 17040 2440
rect 16531 2400 17040 2428
rect 16531 2397 16543 2400
rect 16485 2391 16543 2397
rect 17034 2388 17040 2400
rect 17092 2388 17098 2440
rect 4614 2320 4620 2372
rect 4672 2320 4678 2372
rect 8202 2320 8208 2372
rect 8260 2320 8266 2372
rect 1104 2202 17112 2224
rect 1104 2150 7214 2202
rect 7266 2150 7278 2202
rect 7330 2150 7342 2202
rect 7394 2150 7406 2202
rect 7458 2150 7470 2202
rect 7522 2150 13214 2202
rect 13266 2150 13278 2202
rect 13330 2150 13342 2202
rect 13394 2150 13406 2202
rect 13458 2150 13470 2202
rect 13522 2150 17112 2202
rect 1104 2128 17112 2150
<< via1 >>
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 10214 17926 10266 17978
rect 10278 17926 10330 17978
rect 10342 17926 10394 17978
rect 10406 17926 10458 17978
rect 10470 17926 10522 17978
rect 16214 17926 16266 17978
rect 16278 17926 16330 17978
rect 16342 17926 16394 17978
rect 16406 17926 16458 17978
rect 16470 17926 16522 17978
rect 664 17688 716 17740
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 17040 17688 17092 17740
rect 16212 17620 16264 17672
rect 1584 17527 1636 17536
rect 1584 17493 1593 17527
rect 1593 17493 1627 17527
rect 1627 17493 1636 17527
rect 1584 17484 1636 17493
rect 2688 17527 2740 17536
rect 2688 17493 2697 17527
rect 2697 17493 2731 17527
rect 2731 17493 2740 17527
rect 2688 17484 2740 17493
rect 15936 17527 15988 17536
rect 15936 17493 15945 17527
rect 15945 17493 15979 17527
rect 15979 17493 15988 17527
rect 15936 17484 15988 17493
rect 16212 17527 16264 17536
rect 16212 17493 16221 17527
rect 16221 17493 16255 17527
rect 16255 17493 16264 17527
rect 16212 17484 16264 17493
rect 7214 17382 7266 17434
rect 7278 17382 7330 17434
rect 7342 17382 7394 17434
rect 7406 17382 7458 17434
rect 7470 17382 7522 17434
rect 13214 17382 13266 17434
rect 13278 17382 13330 17434
rect 13342 17382 13394 17434
rect 13406 17382 13458 17434
rect 13470 17382 13522 17434
rect 2596 17280 2648 17332
rect 15936 17280 15988 17332
rect 16212 17280 16264 17332
rect 1584 17144 1636 17196
rect 2044 17144 2096 17196
rect 5448 17144 5500 17196
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 12900 17144 12952 17196
rect 4068 16940 4120 16992
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 11244 16983 11296 16992
rect 11244 16949 11253 16983
rect 11253 16949 11287 16983
rect 11287 16949 11296 16983
rect 11244 16940 11296 16949
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 11888 17076 11940 17128
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 12532 16940 12584 16992
rect 13268 16983 13320 16992
rect 13268 16949 13277 16983
rect 13277 16949 13311 16983
rect 13311 16949 13320 16983
rect 13268 16940 13320 16949
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 10214 16838 10266 16890
rect 10278 16838 10330 16890
rect 10342 16838 10394 16890
rect 10406 16838 10458 16890
rect 10470 16838 10522 16890
rect 16214 16838 16266 16890
rect 16278 16838 16330 16890
rect 16342 16838 16394 16890
rect 16406 16838 16458 16890
rect 16470 16838 16522 16890
rect 2872 16736 2924 16788
rect 11244 16736 11296 16788
rect 11796 16736 11848 16788
rect 13268 16736 13320 16788
rect 2596 16711 2648 16720
rect 2596 16677 2605 16711
rect 2605 16677 2639 16711
rect 2639 16677 2648 16711
rect 2596 16668 2648 16677
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 2136 16532 2188 16584
rect 5540 16532 5592 16584
rect 11428 16532 11480 16584
rect 2320 16507 2372 16516
rect 2320 16473 2329 16507
rect 2329 16473 2363 16507
rect 2363 16473 2372 16507
rect 2320 16464 2372 16473
rect 5448 16464 5500 16516
rect 5540 16439 5592 16448
rect 5540 16405 5549 16439
rect 5549 16405 5583 16439
rect 5583 16405 5592 16439
rect 5540 16396 5592 16405
rect 5816 16439 5868 16448
rect 5816 16405 5825 16439
rect 5825 16405 5859 16439
rect 5859 16405 5868 16439
rect 5816 16396 5868 16405
rect 13820 16532 13872 16584
rect 14188 16575 14240 16584
rect 14188 16541 14197 16575
rect 14197 16541 14231 16575
rect 14231 16541 14240 16575
rect 14188 16532 14240 16541
rect 13268 16464 13320 16516
rect 14556 16464 14608 16516
rect 12624 16396 12676 16448
rect 12716 16396 12768 16448
rect 13360 16396 13412 16448
rect 13544 16439 13596 16448
rect 13544 16405 13553 16439
rect 13553 16405 13587 16439
rect 13587 16405 13596 16439
rect 13544 16396 13596 16405
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 7214 16294 7266 16346
rect 7278 16294 7330 16346
rect 7342 16294 7394 16346
rect 7406 16294 7458 16346
rect 7470 16294 7522 16346
rect 13214 16294 13266 16346
rect 13278 16294 13330 16346
rect 13342 16294 13394 16346
rect 13406 16294 13458 16346
rect 13470 16294 13522 16346
rect 2228 16192 2280 16244
rect 940 16056 992 16108
rect 2136 16056 2188 16108
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 2320 16056 2372 16108
rect 2688 16099 2740 16108
rect 2688 16065 2697 16099
rect 2697 16065 2731 16099
rect 2731 16065 2740 16099
rect 2688 16056 2740 16065
rect 5540 16192 5592 16244
rect 5816 16056 5868 16108
rect 12624 16056 12676 16108
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 13544 16167 13596 16176
rect 13544 16133 13553 16167
rect 13553 16133 13587 16167
rect 13587 16133 13596 16167
rect 13544 16124 13596 16133
rect 14556 16056 14608 16108
rect 14188 15988 14240 16040
rect 2780 15920 2832 15972
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 1768 15852 1820 15904
rect 2688 15895 2740 15904
rect 2688 15861 2697 15895
rect 2697 15861 2731 15895
rect 2731 15861 2740 15895
rect 2688 15852 2740 15861
rect 5264 15895 5316 15904
rect 5264 15861 5273 15895
rect 5273 15861 5307 15895
rect 5307 15861 5316 15895
rect 5264 15852 5316 15861
rect 12532 15895 12584 15904
rect 12532 15861 12541 15895
rect 12541 15861 12575 15895
rect 12575 15861 12584 15895
rect 12532 15852 12584 15861
rect 15476 15852 15528 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 10214 15750 10266 15802
rect 10278 15750 10330 15802
rect 10342 15750 10394 15802
rect 10406 15750 10458 15802
rect 10470 15750 10522 15802
rect 16214 15750 16266 15802
rect 16278 15750 16330 15802
rect 16342 15750 16394 15802
rect 16406 15750 16458 15802
rect 16470 15750 16522 15802
rect 13084 15648 13136 15700
rect 14280 15648 14332 15700
rect 5448 15580 5500 15632
rect 1768 15555 1820 15564
rect 1768 15521 1777 15555
rect 1777 15521 1811 15555
rect 1811 15521 1820 15555
rect 1768 15512 1820 15521
rect 2688 15512 2740 15564
rect 11428 15580 11480 15632
rect 5356 15444 5408 15496
rect 4160 15376 4212 15428
rect 6092 15376 6144 15428
rect 9036 15444 9088 15496
rect 15476 15512 15528 15564
rect 8300 15376 8352 15428
rect 8668 15376 8720 15428
rect 10968 15376 11020 15428
rect 14372 15376 14424 15428
rect 14556 15376 14608 15428
rect 3332 15308 3384 15360
rect 4804 15351 4856 15360
rect 4804 15317 4813 15351
rect 4813 15317 4847 15351
rect 4847 15317 4856 15351
rect 4804 15308 4856 15317
rect 7104 15308 7156 15360
rect 8484 15351 8536 15360
rect 8484 15317 8493 15351
rect 8493 15317 8527 15351
rect 8527 15317 8536 15351
rect 8484 15308 8536 15317
rect 9312 15308 9364 15360
rect 11336 15308 11388 15360
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 7214 15206 7266 15258
rect 7278 15206 7330 15258
rect 7342 15206 7394 15258
rect 7406 15206 7458 15258
rect 7470 15206 7522 15258
rect 13214 15206 13266 15258
rect 13278 15206 13330 15258
rect 13342 15206 13394 15258
rect 13406 15206 13458 15258
rect 13470 15206 13522 15258
rect 5356 15147 5408 15156
rect 5356 15113 5365 15147
rect 5365 15113 5399 15147
rect 5399 15113 5408 15147
rect 5356 15104 5408 15113
rect 8668 15147 8720 15156
rect 8668 15113 8677 15147
rect 8677 15113 8711 15147
rect 8711 15113 8720 15147
rect 8668 15104 8720 15113
rect 9036 15104 9088 15156
rect 10692 15104 10744 15156
rect 1768 15036 1820 15088
rect 3332 15036 3384 15088
rect 7104 15036 7156 15088
rect 8484 15036 8536 15088
rect 14188 15104 14240 15156
rect 10968 15036 11020 15088
rect 13820 15079 13872 15088
rect 13820 15045 13829 15079
rect 13829 15045 13863 15079
rect 13863 15045 13872 15079
rect 13820 15036 13872 15045
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 4160 14968 4212 15020
rect 4620 14968 4672 15020
rect 4804 15011 4856 15020
rect 4804 14977 4813 15011
rect 4813 14977 4847 15011
rect 4847 14977 4856 15011
rect 4804 14968 4856 14977
rect 5264 14968 5316 15020
rect 6092 14968 6144 15020
rect 6828 14968 6880 15020
rect 8300 14968 8352 15020
rect 8668 14968 8720 15020
rect 8944 14968 8996 15020
rect 9036 15011 9088 15020
rect 9036 14977 9045 15011
rect 9045 14977 9079 15011
rect 9079 14977 9088 15011
rect 9036 14968 9088 14977
rect 2228 14900 2280 14952
rect 9588 14968 9640 15020
rect 11428 14968 11480 15020
rect 11612 14968 11664 15020
rect 11060 14943 11112 14952
rect 11060 14909 11069 14943
rect 11069 14909 11103 14943
rect 11103 14909 11112 14943
rect 11060 14900 11112 14909
rect 11336 14943 11388 14952
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 9680 14832 9732 14884
rect 15936 14968 15988 15020
rect 15292 14943 15344 14952
rect 15292 14909 15301 14943
rect 15301 14909 15335 14943
rect 15335 14909 15344 14943
rect 15292 14900 15344 14909
rect 2504 14807 2556 14816
rect 2504 14773 2513 14807
rect 2513 14773 2547 14807
rect 2547 14773 2556 14807
rect 2504 14764 2556 14773
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 9404 14764 9456 14773
rect 12440 14764 12492 14816
rect 12808 14764 12860 14816
rect 12992 14764 13044 14816
rect 13544 14764 13596 14816
rect 15568 14764 15620 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 10214 14662 10266 14714
rect 10278 14662 10330 14714
rect 10342 14662 10394 14714
rect 10406 14662 10458 14714
rect 10470 14662 10522 14714
rect 16214 14662 16266 14714
rect 16278 14662 16330 14714
rect 16342 14662 16394 14714
rect 16406 14662 16458 14714
rect 16470 14662 16522 14714
rect 4804 14560 4856 14612
rect 6828 14560 6880 14612
rect 8484 14560 8536 14612
rect 11060 14560 11112 14612
rect 11428 14560 11480 14612
rect 12256 14603 12308 14612
rect 12256 14569 12265 14603
rect 12265 14569 12299 14603
rect 12299 14569 12308 14603
rect 12256 14560 12308 14569
rect 13820 14603 13872 14612
rect 13820 14569 13829 14603
rect 13829 14569 13863 14603
rect 13863 14569 13872 14603
rect 13820 14560 13872 14569
rect 15936 14560 15988 14612
rect 9312 14424 9364 14476
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 10968 14356 11020 14408
rect 11612 14424 11664 14476
rect 12440 14492 12492 14544
rect 12256 14356 12308 14408
rect 7840 14288 7892 14340
rect 3976 14263 4028 14272
rect 3976 14229 3985 14263
rect 3985 14229 4019 14263
rect 4019 14229 4028 14263
rect 3976 14220 4028 14229
rect 10692 14288 10744 14340
rect 13084 14288 13136 14340
rect 14280 14220 14332 14272
rect 15568 14399 15620 14408
rect 15568 14365 15602 14399
rect 15602 14365 15620 14399
rect 15568 14356 15620 14365
rect 7214 14118 7266 14170
rect 7278 14118 7330 14170
rect 7342 14118 7394 14170
rect 7406 14118 7458 14170
rect 7470 14118 7522 14170
rect 13214 14118 13266 14170
rect 13278 14118 13330 14170
rect 13342 14118 13394 14170
rect 13406 14118 13458 14170
rect 13470 14118 13522 14170
rect 3976 14016 4028 14068
rect 7840 14059 7892 14068
rect 7840 14025 7849 14059
rect 7849 14025 7883 14059
rect 7883 14025 7892 14059
rect 7840 14016 7892 14025
rect 8944 14016 8996 14068
rect 13084 14059 13136 14068
rect 13084 14025 13093 14059
rect 13093 14025 13127 14059
rect 13127 14025 13136 14059
rect 13084 14016 13136 14025
rect 13544 14016 13596 14068
rect 15476 14016 15528 14068
rect 9404 13948 9456 14000
rect 12992 13923 13044 13932
rect 12992 13889 13001 13923
rect 13001 13889 13035 13923
rect 13035 13889 13044 13923
rect 12992 13880 13044 13889
rect 14648 13880 14700 13932
rect 16028 13880 16080 13932
rect 10140 13855 10192 13864
rect 10140 13821 10149 13855
rect 10149 13821 10183 13855
rect 10183 13821 10192 13855
rect 10140 13812 10192 13821
rect 12256 13812 12308 13864
rect 3424 13719 3476 13728
rect 3424 13685 3433 13719
rect 3433 13685 3467 13719
rect 3467 13685 3476 13719
rect 3424 13676 3476 13685
rect 14280 13676 14332 13728
rect 15568 13719 15620 13728
rect 15568 13685 15577 13719
rect 15577 13685 15611 13719
rect 15611 13685 15620 13719
rect 15568 13676 15620 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 10214 13574 10266 13626
rect 10278 13574 10330 13626
rect 10342 13574 10394 13626
rect 10406 13574 10458 13626
rect 10470 13574 10522 13626
rect 16214 13574 16266 13626
rect 16278 13574 16330 13626
rect 16342 13574 16394 13626
rect 16406 13574 16458 13626
rect 16470 13574 16522 13626
rect 14648 13515 14700 13524
rect 14648 13481 14657 13515
rect 14657 13481 14691 13515
rect 14691 13481 14700 13515
rect 14648 13472 14700 13481
rect 15292 13472 15344 13524
rect 9404 13336 9456 13388
rect 10416 13336 10468 13388
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 6276 13311 6328 13320
rect 6276 13277 6285 13311
rect 6285 13277 6319 13311
rect 6319 13277 6328 13311
rect 6276 13268 6328 13277
rect 10692 13268 10744 13320
rect 12440 13268 12492 13320
rect 13820 13311 13872 13320
rect 13820 13277 13829 13311
rect 13829 13277 13863 13311
rect 13863 13277 13872 13311
rect 13820 13268 13872 13277
rect 6552 13243 6604 13252
rect 6552 13209 6561 13243
rect 6561 13209 6595 13243
rect 6595 13209 6604 13243
rect 6552 13200 6604 13209
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 4620 13132 4672 13184
rect 8300 13200 8352 13252
rect 8852 13200 8904 13252
rect 9312 13200 9364 13252
rect 13544 13243 13596 13252
rect 13544 13209 13553 13243
rect 13553 13209 13587 13243
rect 13587 13209 13596 13243
rect 13544 13200 13596 13209
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 15568 13268 15620 13320
rect 8024 13175 8076 13184
rect 8024 13141 8033 13175
rect 8033 13141 8067 13175
rect 8067 13141 8076 13175
rect 8024 13132 8076 13141
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 16028 13132 16080 13184
rect 7214 13030 7266 13082
rect 7278 13030 7330 13082
rect 7342 13030 7394 13082
rect 7406 13030 7458 13082
rect 7470 13030 7522 13082
rect 13214 13030 13266 13082
rect 13278 13030 13330 13082
rect 13342 13030 13394 13082
rect 13406 13030 13458 13082
rect 13470 13030 13522 13082
rect 2504 12860 2556 12912
rect 4896 12792 4948 12844
rect 6276 12792 6328 12844
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 6920 12767 6972 12776
rect 6920 12733 6929 12767
rect 6929 12733 6963 12767
rect 6963 12733 6972 12767
rect 6920 12724 6972 12733
rect 7104 12835 7156 12844
rect 7104 12801 7113 12835
rect 7113 12801 7147 12835
rect 7147 12801 7156 12835
rect 7104 12792 7156 12801
rect 8024 12928 8076 12980
rect 9312 12971 9364 12980
rect 9312 12937 9321 12971
rect 9321 12937 9355 12971
rect 9355 12937 9364 12971
rect 9312 12928 9364 12937
rect 8300 12860 8352 12912
rect 10600 12928 10652 12980
rect 10784 12928 10836 12980
rect 13544 12928 13596 12980
rect 9496 12792 9548 12844
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 5264 12699 5316 12708
rect 5264 12665 5273 12699
rect 5273 12665 5307 12699
rect 5307 12665 5316 12699
rect 5264 12656 5316 12665
rect 5908 12656 5960 12708
rect 6644 12699 6696 12708
rect 6644 12665 6653 12699
rect 6653 12665 6687 12699
rect 6687 12665 6696 12699
rect 6644 12656 6696 12665
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 6460 12631 6512 12640
rect 6460 12597 6469 12631
rect 6469 12597 6503 12631
rect 6503 12597 6512 12631
rect 6460 12588 6512 12597
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 10416 12792 10468 12844
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 12440 12860 12492 12912
rect 15016 12860 15068 12912
rect 15200 12860 15252 12912
rect 15844 12792 15896 12844
rect 9864 12588 9916 12640
rect 12532 12724 12584 12776
rect 10600 12699 10652 12708
rect 10600 12665 10609 12699
rect 10609 12665 10643 12699
rect 10643 12665 10652 12699
rect 10600 12656 10652 12665
rect 12256 12588 12308 12640
rect 14280 12631 14332 12640
rect 14280 12597 14289 12631
rect 14289 12597 14323 12631
rect 14323 12597 14332 12631
rect 14280 12588 14332 12597
rect 15292 12631 15344 12640
rect 15292 12597 15301 12631
rect 15301 12597 15335 12631
rect 15335 12597 15344 12631
rect 15292 12588 15344 12597
rect 16028 12588 16080 12640
rect 16120 12588 16172 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 10214 12486 10266 12538
rect 10278 12486 10330 12538
rect 10342 12486 10394 12538
rect 10406 12486 10458 12538
rect 10470 12486 10522 12538
rect 16214 12486 16266 12538
rect 16278 12486 16330 12538
rect 16342 12486 16394 12538
rect 16406 12486 16458 12538
rect 16470 12486 16522 12538
rect 6552 12384 6604 12436
rect 12256 12427 12308 12436
rect 12256 12393 12265 12427
rect 12265 12393 12299 12427
rect 12299 12393 12308 12427
rect 12256 12384 12308 12393
rect 13820 12384 13872 12436
rect 6276 12316 6328 12368
rect 7104 12316 7156 12368
rect 12532 12316 12584 12368
rect 13084 12316 13136 12368
rect 1676 12248 1728 12300
rect 10140 12248 10192 12300
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 5264 12180 5316 12232
rect 6460 12180 6512 12232
rect 14924 12248 14976 12300
rect 2136 12155 2188 12164
rect 2136 12121 2145 12155
rect 2145 12121 2179 12155
rect 2179 12121 2188 12155
rect 2136 12112 2188 12121
rect 3700 12112 3752 12164
rect 4620 12112 4672 12164
rect 12440 12112 12492 12164
rect 3424 12044 3476 12096
rect 12716 12044 12768 12096
rect 14280 12180 14332 12232
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 13728 12155 13780 12164
rect 13728 12121 13737 12155
rect 13737 12121 13771 12155
rect 13771 12121 13780 12155
rect 13728 12112 13780 12121
rect 14188 12044 14240 12096
rect 15292 12112 15344 12164
rect 7214 11942 7266 11994
rect 7278 11942 7330 11994
rect 7342 11942 7394 11994
rect 7406 11942 7458 11994
rect 7470 11942 7522 11994
rect 13214 11942 13266 11994
rect 13278 11942 13330 11994
rect 13342 11942 13394 11994
rect 13406 11942 13458 11994
rect 13470 11942 13522 11994
rect 3424 11840 3476 11892
rect 4712 11840 4764 11892
rect 6920 11840 6972 11892
rect 4620 11772 4672 11824
rect 7104 11772 7156 11824
rect 2872 11747 2924 11756
rect 2872 11713 2881 11747
rect 2881 11713 2915 11747
rect 2915 11713 2924 11747
rect 2872 11704 2924 11713
rect 4160 11568 4212 11620
rect 4804 11704 4856 11756
rect 4896 11747 4948 11756
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 6644 11704 6696 11756
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 9128 11704 9180 11756
rect 9680 11815 9732 11824
rect 9680 11781 9689 11815
rect 9689 11781 9723 11815
rect 9723 11781 9732 11815
rect 9680 11772 9732 11781
rect 9864 11704 9916 11756
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 12808 11704 12860 11756
rect 13084 11840 13136 11892
rect 14188 11840 14240 11892
rect 15108 11840 15160 11892
rect 14280 11772 14332 11824
rect 13544 11704 13596 11756
rect 15292 11747 15344 11756
rect 15292 11713 15326 11747
rect 15326 11713 15344 11747
rect 15292 11704 15344 11713
rect 11152 11568 11204 11620
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 7932 11543 7984 11552
rect 7932 11509 7941 11543
rect 7941 11509 7975 11543
rect 7975 11509 7984 11543
rect 7932 11500 7984 11509
rect 8852 11500 8904 11552
rect 11336 11500 11388 11552
rect 11428 11500 11480 11552
rect 13268 11500 13320 11552
rect 15016 11500 15068 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 10214 11398 10266 11450
rect 10278 11398 10330 11450
rect 10342 11398 10394 11450
rect 10406 11398 10458 11450
rect 10470 11398 10522 11450
rect 16214 11398 16266 11450
rect 16278 11398 16330 11450
rect 16342 11398 16394 11450
rect 16406 11398 16458 11450
rect 16470 11398 16522 11450
rect 2136 11296 2188 11348
rect 7012 11296 7064 11348
rect 7932 11296 7984 11348
rect 4620 11271 4672 11280
rect 4620 11237 4629 11271
rect 4629 11237 4663 11271
rect 4663 11237 4672 11271
rect 4620 11228 4672 11237
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 5724 11160 5776 11212
rect 11152 11296 11204 11348
rect 11336 11296 11388 11348
rect 13268 11296 13320 11348
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 15292 11296 15344 11348
rect 4804 11092 4856 11144
rect 4988 11092 5040 11144
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 4344 11067 4396 11076
rect 4344 11033 4353 11067
rect 4353 11033 4387 11067
rect 4387 11033 4396 11067
rect 4344 11024 4396 11033
rect 6828 11092 6880 11144
rect 12440 11160 12492 11212
rect 13084 11092 13136 11144
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 15200 11160 15252 11212
rect 13728 11092 13780 11101
rect 8852 11024 8904 11076
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 12440 11024 12492 11076
rect 15016 11024 15068 11076
rect 4712 10956 4764 11008
rect 4896 10956 4948 11008
rect 5816 10999 5868 11008
rect 5816 10965 5825 10999
rect 5825 10965 5859 10999
rect 5859 10965 5868 10999
rect 5816 10956 5868 10965
rect 6276 10956 6328 11008
rect 8668 10999 8720 11008
rect 8668 10965 8677 10999
rect 8677 10965 8711 10999
rect 8711 10965 8720 10999
rect 8668 10956 8720 10965
rect 12624 10956 12676 11008
rect 7214 10854 7266 10906
rect 7278 10854 7330 10906
rect 7342 10854 7394 10906
rect 7406 10854 7458 10906
rect 7470 10854 7522 10906
rect 13214 10854 13266 10906
rect 13278 10854 13330 10906
rect 13342 10854 13394 10906
rect 13406 10854 13458 10906
rect 13470 10854 13522 10906
rect 4344 10752 4396 10804
rect 4804 10752 4856 10804
rect 6000 10752 6052 10804
rect 7656 10752 7708 10804
rect 9864 10795 9916 10804
rect 9864 10761 9873 10795
rect 9873 10761 9907 10795
rect 9907 10761 9916 10795
rect 9864 10752 9916 10761
rect 10140 10752 10192 10804
rect 2780 10659 2832 10668
rect 2780 10625 2789 10659
rect 2789 10625 2823 10659
rect 2823 10625 2832 10659
rect 2780 10616 2832 10625
rect 940 10548 992 10600
rect 4620 10616 4672 10668
rect 5540 10616 5592 10668
rect 6276 10616 6328 10668
rect 4712 10548 4764 10600
rect 6828 10684 6880 10736
rect 8668 10684 8720 10736
rect 8852 10684 8904 10736
rect 12256 10684 12308 10736
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15200 10659 15252 10668
rect 15200 10625 15214 10659
rect 15214 10625 15248 10659
rect 15248 10625 15252 10659
rect 15200 10616 15252 10625
rect 15476 10616 15528 10668
rect 11244 10591 11296 10600
rect 11244 10557 11253 10591
rect 11253 10557 11287 10591
rect 11287 10557 11296 10591
rect 11244 10548 11296 10557
rect 13084 10548 13136 10600
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 15844 10548 15896 10600
rect 3332 10455 3384 10464
rect 3332 10421 3341 10455
rect 3341 10421 3375 10455
rect 3375 10421 3384 10455
rect 3332 10412 3384 10421
rect 11520 10412 11572 10464
rect 13360 10455 13412 10464
rect 13360 10421 13369 10455
rect 13369 10421 13403 10455
rect 13403 10421 13412 10455
rect 13360 10412 13412 10421
rect 14188 10455 14240 10464
rect 14188 10421 14197 10455
rect 14197 10421 14231 10455
rect 14231 10421 14240 10455
rect 14188 10412 14240 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 10214 10310 10266 10362
rect 10278 10310 10330 10362
rect 10342 10310 10394 10362
rect 10406 10310 10458 10362
rect 10470 10310 10522 10362
rect 16214 10310 16266 10362
rect 16278 10310 16330 10362
rect 16342 10310 16394 10362
rect 16406 10310 16458 10362
rect 16470 10310 16522 10362
rect 3056 10208 3108 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 2872 10140 2924 10192
rect 4620 10183 4672 10192
rect 4620 10149 4629 10183
rect 4629 10149 4663 10183
rect 4663 10149 4672 10183
rect 4620 10140 4672 10149
rect 4068 10047 4120 10056
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4804 10004 4856 10056
rect 4988 10004 5040 10056
rect 5816 10004 5868 10056
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 6368 10047 6420 10056
rect 6368 10013 6377 10047
rect 6377 10013 6411 10047
rect 6411 10013 6420 10047
rect 6368 10004 6420 10013
rect 11244 10140 11296 10192
rect 11336 10183 11388 10192
rect 11336 10149 11345 10183
rect 11345 10149 11379 10183
rect 11379 10149 11388 10183
rect 11336 10140 11388 10149
rect 12624 10208 12676 10260
rect 12900 10208 12952 10260
rect 14372 10208 14424 10260
rect 11152 10047 11204 10056
rect 11152 10013 11166 10047
rect 11166 10013 11200 10047
rect 11200 10013 11204 10047
rect 11152 10004 11204 10013
rect 11520 10047 11572 10056
rect 11520 10013 11529 10047
rect 11529 10013 11563 10047
rect 11563 10013 11572 10047
rect 11520 10004 11572 10013
rect 12256 10072 12308 10124
rect 16120 10072 16172 10124
rect 13360 10004 13412 10056
rect 3148 9868 3200 9920
rect 3700 9868 3752 9920
rect 10968 9979 11020 9988
rect 10968 9945 10977 9979
rect 10977 9945 11011 9979
rect 11011 9945 11020 9979
rect 10968 9936 11020 9945
rect 4436 9868 4488 9920
rect 4528 9868 4580 9920
rect 6276 9868 6328 9920
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 11152 9868 11204 9920
rect 12532 9936 12584 9988
rect 14740 10004 14792 10056
rect 13912 9936 13964 9988
rect 15752 9936 15804 9988
rect 13636 9868 13688 9920
rect 14464 9868 14516 9920
rect 15108 9868 15160 9920
rect 15844 9868 15896 9920
rect 7214 9766 7266 9818
rect 7278 9766 7330 9818
rect 7342 9766 7394 9818
rect 7406 9766 7458 9818
rect 7470 9766 7522 9818
rect 13214 9766 13266 9818
rect 13278 9766 13330 9818
rect 13342 9766 13394 9818
rect 13406 9766 13458 9818
rect 13470 9766 13522 9818
rect 1860 9664 1912 9716
rect 2780 9664 2832 9716
rect 3056 9664 3108 9716
rect 4528 9707 4580 9716
rect 4528 9673 4537 9707
rect 4537 9673 4571 9707
rect 4571 9673 4580 9707
rect 4528 9664 4580 9673
rect 4620 9664 4672 9716
rect 11244 9707 11296 9716
rect 11244 9673 11253 9707
rect 11253 9673 11287 9707
rect 11287 9673 11296 9707
rect 11244 9664 11296 9673
rect 11336 9664 11388 9716
rect 12256 9664 12308 9716
rect 12532 9664 12584 9716
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 3700 9596 3752 9648
rect 8576 9596 8628 9648
rect 10876 9528 10928 9580
rect 14188 9664 14240 9716
rect 14832 9664 14884 9716
rect 3148 9460 3200 9512
rect 4896 9324 4948 9376
rect 6460 9324 6512 9376
rect 7656 9324 7708 9376
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 11152 9324 11204 9376
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 14004 9596 14056 9648
rect 15844 9664 15896 9716
rect 13544 9460 13596 9512
rect 15476 9571 15528 9580
rect 15476 9537 15477 9571
rect 15477 9537 15511 9571
rect 15511 9537 15528 9571
rect 15476 9528 15528 9537
rect 14464 9324 14516 9376
rect 15016 9367 15068 9376
rect 15016 9333 15025 9367
rect 15025 9333 15059 9367
rect 15059 9333 15068 9367
rect 15016 9324 15068 9333
rect 15384 9324 15436 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 10214 9222 10266 9274
rect 10278 9222 10330 9274
rect 10342 9222 10394 9274
rect 10406 9222 10458 9274
rect 10470 9222 10522 9274
rect 16214 9222 16266 9274
rect 16278 9222 16330 9274
rect 16342 9222 16394 9274
rect 16406 9222 16458 9274
rect 16470 9222 16522 9274
rect 2412 9120 2464 9172
rect 6276 9052 6328 9104
rect 6460 8984 6512 9036
rect 1860 8916 1912 8968
rect 6092 8916 6144 8968
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 11428 9163 11480 9172
rect 11428 9129 11437 9163
rect 11437 9129 11471 9163
rect 11471 9129 11480 9163
rect 11428 9120 11480 9129
rect 13912 9163 13964 9172
rect 13912 9129 13921 9163
rect 13921 9129 13955 9163
rect 13955 9129 13964 9163
rect 13912 9120 13964 9129
rect 7656 9052 7708 9104
rect 4896 8848 4948 8900
rect 4988 8891 5040 8900
rect 4988 8857 4997 8891
rect 4997 8857 5031 8891
rect 5031 8857 5040 8891
rect 4988 8848 5040 8857
rect 1584 8780 1636 8832
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 7748 8984 7800 9036
rect 13636 8984 13688 9036
rect 15016 8984 15068 9036
rect 16120 9163 16172 9172
rect 16120 9129 16129 9163
rect 16129 9129 16163 9163
rect 16163 9129 16172 9163
rect 16120 9120 16172 9129
rect 10968 8916 11020 8968
rect 6460 8780 6512 8789
rect 7564 8780 7616 8832
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 13084 8848 13136 8900
rect 13544 8780 13596 8832
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 15752 8916 15804 8968
rect 15384 8780 15436 8832
rect 7214 8678 7266 8730
rect 7278 8678 7330 8730
rect 7342 8678 7394 8730
rect 7406 8678 7458 8730
rect 7470 8678 7522 8730
rect 13214 8678 13266 8730
rect 13278 8678 13330 8730
rect 13342 8678 13394 8730
rect 13406 8678 13458 8730
rect 13470 8678 13522 8730
rect 4988 8576 5040 8628
rect 7748 8576 7800 8628
rect 13084 8576 13136 8628
rect 13544 8576 13596 8628
rect 14372 8576 14424 8628
rect 15476 8576 15528 8628
rect 6092 8508 6144 8560
rect 6460 8508 6512 8560
rect 3332 8440 3384 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 8392 8508 8444 8560
rect 8576 8508 8628 8560
rect 10876 8440 10928 8492
rect 11428 8440 11480 8492
rect 11612 8440 11664 8492
rect 7564 8372 7616 8424
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 13820 8440 13872 8492
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 15108 8440 15160 8492
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 5816 8304 5868 8356
rect 11244 8304 11296 8356
rect 15476 8372 15528 8424
rect 13360 8347 13412 8356
rect 13360 8313 13369 8347
rect 13369 8313 13403 8347
rect 13403 8313 13412 8347
rect 13360 8304 13412 8313
rect 6920 8279 6972 8288
rect 6920 8245 6929 8279
rect 6929 8245 6963 8279
rect 6963 8245 6972 8279
rect 6920 8236 6972 8245
rect 14556 8279 14608 8288
rect 14556 8245 14565 8279
rect 14565 8245 14599 8279
rect 14599 8245 14608 8279
rect 14556 8236 14608 8245
rect 14740 8279 14792 8288
rect 14740 8245 14749 8279
rect 14749 8245 14783 8279
rect 14783 8245 14792 8279
rect 14740 8236 14792 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 10214 8134 10266 8186
rect 10278 8134 10330 8186
rect 10342 8134 10394 8186
rect 10406 8134 10458 8186
rect 10470 8134 10522 8186
rect 16214 8134 16266 8186
rect 16278 8134 16330 8186
rect 16342 8134 16394 8186
rect 16406 8134 16458 8186
rect 16470 8134 16522 8186
rect 8392 8075 8444 8084
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 11612 8075 11664 8084
rect 11612 8041 11621 8075
rect 11621 8041 11655 8075
rect 11655 8041 11664 8075
rect 11612 8032 11664 8041
rect 13636 8032 13688 8084
rect 6276 7896 6328 7948
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 9588 7828 9640 7880
rect 11244 7828 11296 7880
rect 14740 8032 14792 8084
rect 14372 7896 14424 7948
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 8576 7760 8628 7812
rect 9772 7803 9824 7812
rect 9772 7769 9806 7803
rect 9806 7769 9824 7803
rect 9772 7760 9824 7769
rect 15108 7760 15160 7812
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 2780 7692 2832 7701
rect 6092 7692 6144 7744
rect 8208 7692 8260 7744
rect 15844 7735 15896 7744
rect 15844 7701 15853 7735
rect 15853 7701 15887 7735
rect 15887 7701 15896 7735
rect 15844 7692 15896 7701
rect 7214 7590 7266 7642
rect 7278 7590 7330 7642
rect 7342 7590 7394 7642
rect 7406 7590 7458 7642
rect 7470 7590 7522 7642
rect 13214 7590 13266 7642
rect 13278 7590 13330 7642
rect 13342 7590 13394 7642
rect 13406 7590 13458 7642
rect 13470 7590 13522 7642
rect 2780 7488 2832 7540
rect 4620 7488 4672 7540
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 11428 7488 11480 7540
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 15476 7488 15528 7540
rect 15844 7488 15896 7540
rect 6092 7420 6144 7472
rect 9496 7395 9548 7404
rect 9496 7361 9505 7395
rect 9505 7361 9539 7395
rect 9539 7361 9548 7395
rect 9496 7352 9548 7361
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 10968 7420 11020 7472
rect 12716 7420 12768 7472
rect 14556 7420 14608 7472
rect 11428 7352 11480 7404
rect 15108 7352 15160 7404
rect 16580 7352 16632 7404
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 16580 7216 16632 7268
rect 4620 7148 4672 7200
rect 6000 7148 6052 7200
rect 12992 7148 13044 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 10214 7046 10266 7098
rect 10278 7046 10330 7098
rect 10342 7046 10394 7098
rect 10406 7046 10458 7098
rect 10470 7046 10522 7098
rect 16214 7046 16266 7098
rect 16278 7046 16330 7098
rect 16342 7046 16394 7098
rect 16406 7046 16458 7098
rect 16470 7046 16522 7098
rect 6000 6987 6052 6996
rect 6000 6953 6030 6987
rect 6030 6953 6052 6987
rect 6000 6944 6052 6953
rect 7656 6808 7708 6860
rect 8116 6808 8168 6860
rect 9588 6944 9640 6996
rect 9680 6876 9732 6928
rect 12716 6944 12768 6996
rect 13636 6944 13688 6996
rect 16580 6987 16632 6996
rect 16580 6953 16589 6987
rect 16589 6953 16623 6987
rect 16623 6953 16632 6987
rect 16580 6944 16632 6953
rect 11428 6876 11480 6928
rect 8760 6740 8812 6792
rect 8208 6672 8260 6724
rect 7012 6604 7064 6656
rect 8024 6604 8076 6656
rect 8116 6604 8168 6656
rect 10140 6851 10192 6860
rect 10140 6817 10149 6851
rect 10149 6817 10183 6851
rect 10183 6817 10192 6851
rect 10140 6808 10192 6817
rect 12072 6808 12124 6860
rect 12348 6851 12400 6860
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 12440 6851 12492 6860
rect 12440 6817 12450 6851
rect 12450 6817 12484 6851
rect 12484 6817 12492 6851
rect 12440 6808 12492 6817
rect 12900 6919 12952 6928
rect 12900 6885 12909 6919
rect 12909 6885 12943 6919
rect 12943 6885 12952 6919
rect 12900 6876 12952 6885
rect 17132 6808 17184 6860
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 9956 6604 10008 6656
rect 10416 6715 10468 6724
rect 10416 6681 10425 6715
rect 10425 6681 10459 6715
rect 10459 6681 10468 6715
rect 10416 6672 10468 6681
rect 10968 6672 11020 6724
rect 13728 6740 13780 6792
rect 10784 6604 10836 6656
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 12348 6604 12400 6656
rect 12992 6672 13044 6724
rect 7214 6502 7266 6554
rect 7278 6502 7330 6554
rect 7342 6502 7394 6554
rect 7406 6502 7458 6554
rect 7470 6502 7522 6554
rect 13214 6502 13266 6554
rect 13278 6502 13330 6554
rect 13342 6502 13394 6554
rect 13406 6502 13458 6554
rect 13470 6502 13522 6554
rect 8760 6443 8812 6452
rect 8760 6409 8769 6443
rect 8769 6409 8803 6443
rect 8803 6409 8812 6443
rect 8760 6400 8812 6409
rect 10140 6400 10192 6452
rect 10416 6400 10468 6452
rect 11980 6400 12032 6452
rect 12256 6400 12308 6452
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 5172 6332 5224 6384
rect 4620 6264 4672 6273
rect 4988 6307 5040 6316
rect 4988 6273 5022 6307
rect 5022 6273 5040 6307
rect 4988 6264 5040 6273
rect 7012 6264 7064 6316
rect 7840 6332 7892 6384
rect 7656 6307 7708 6316
rect 7656 6273 7690 6307
rect 7690 6273 7708 6307
rect 7656 6264 7708 6273
rect 11152 6264 11204 6316
rect 13912 6400 13964 6452
rect 15660 6400 15712 6452
rect 12900 6264 12952 6316
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 9496 6196 9548 6248
rect 12256 6196 12308 6248
rect 12164 6128 12216 6180
rect 12992 6128 13044 6180
rect 5816 6060 5868 6112
rect 13912 6060 13964 6112
rect 14740 6060 14792 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 10214 5958 10266 6010
rect 10278 5958 10330 6010
rect 10342 5958 10394 6010
rect 10406 5958 10458 6010
rect 10470 5958 10522 6010
rect 16214 5958 16266 6010
rect 16278 5958 16330 6010
rect 16342 5958 16394 6010
rect 16406 5958 16458 6010
rect 16470 5958 16522 6010
rect 2688 5856 2740 5908
rect 4988 5856 5040 5908
rect 5816 5720 5868 5772
rect 4896 5652 4948 5704
rect 8024 5652 8076 5704
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 9956 5695 10008 5704
rect 9956 5661 9965 5695
rect 9965 5661 9999 5695
rect 9999 5661 10008 5695
rect 9956 5652 10008 5661
rect 11152 5899 11204 5908
rect 11152 5865 11161 5899
rect 11161 5865 11195 5899
rect 11195 5865 11204 5899
rect 11152 5856 11204 5865
rect 13636 5856 13688 5908
rect 11888 5720 11940 5772
rect 12532 5720 12584 5772
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 3424 5627 3476 5636
rect 3424 5593 3433 5627
rect 3433 5593 3467 5627
rect 3467 5593 3476 5627
rect 3424 5584 3476 5593
rect 12072 5652 12124 5704
rect 12256 5652 12308 5704
rect 12808 5652 12860 5704
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 7840 5516 7892 5568
rect 9588 5516 9640 5568
rect 10784 5584 10836 5636
rect 12348 5584 12400 5636
rect 13912 5627 13964 5636
rect 13912 5593 13921 5627
rect 13921 5593 13955 5627
rect 13955 5593 13964 5627
rect 13912 5584 13964 5593
rect 15200 5627 15252 5636
rect 15200 5593 15209 5627
rect 15209 5593 15243 5627
rect 15243 5593 15252 5627
rect 15200 5584 15252 5593
rect 15660 5584 15712 5636
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 11612 5559 11664 5568
rect 11612 5525 11621 5559
rect 11621 5525 11655 5559
rect 11655 5525 11664 5559
rect 11612 5516 11664 5525
rect 13820 5516 13872 5568
rect 14740 5516 14792 5568
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 16672 5516 16724 5525
rect 7214 5414 7266 5466
rect 7278 5414 7330 5466
rect 7342 5414 7394 5466
rect 7406 5414 7458 5466
rect 7470 5414 7522 5466
rect 13214 5414 13266 5466
rect 13278 5414 13330 5466
rect 13342 5414 13394 5466
rect 13406 5414 13458 5466
rect 13470 5414 13522 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 4896 5355 4948 5364
rect 4896 5321 4905 5355
rect 4905 5321 4939 5355
rect 4939 5321 4948 5355
rect 4896 5312 4948 5321
rect 11060 5312 11112 5364
rect 5632 5244 5684 5296
rect 940 5176 992 5228
rect 4068 5176 4120 5228
rect 5356 5176 5408 5228
rect 8024 5244 8076 5296
rect 11612 5244 11664 5296
rect 12072 5287 12124 5296
rect 12072 5253 12081 5287
rect 12081 5253 12115 5287
rect 12115 5253 12124 5287
rect 12072 5244 12124 5253
rect 12256 5244 12308 5296
rect 15200 5312 15252 5364
rect 12808 5244 12860 5296
rect 3516 5151 3568 5160
rect 3516 5117 3525 5151
rect 3525 5117 3559 5151
rect 3559 5117 3568 5151
rect 3516 5108 3568 5117
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 8116 5108 8168 5160
rect 8208 5108 8260 5160
rect 7564 5040 7616 5092
rect 5264 4972 5316 5024
rect 5540 4972 5592 5024
rect 5816 4972 5868 5024
rect 6368 4972 6420 5024
rect 6736 4972 6788 5024
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 7196 4972 7248 4981
rect 9772 5108 9824 5160
rect 11244 5108 11296 5160
rect 11520 5083 11572 5092
rect 11520 5049 11529 5083
rect 11529 5049 11563 5083
rect 11563 5049 11572 5083
rect 11520 5040 11572 5049
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 11980 5176 12032 5228
rect 13820 5219 13872 5228
rect 13820 5185 13837 5219
rect 13837 5185 13872 5219
rect 13820 5176 13872 5185
rect 14004 5219 14056 5228
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 14648 5244 14700 5296
rect 16672 5244 16724 5296
rect 14556 5108 14608 5160
rect 12164 4972 12216 5024
rect 12992 4972 13044 5024
rect 13268 4972 13320 5024
rect 14004 4972 14056 5024
rect 14464 4972 14516 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 10214 4870 10266 4922
rect 10278 4870 10330 4922
rect 10342 4870 10394 4922
rect 10406 4870 10458 4922
rect 10470 4870 10522 4922
rect 16214 4870 16266 4922
rect 16278 4870 16330 4922
rect 16342 4870 16394 4922
rect 16406 4870 16458 4922
rect 16470 4870 16522 4922
rect 4068 4768 4120 4820
rect 5632 4768 5684 4820
rect 7012 4768 7064 4820
rect 8208 4768 8260 4820
rect 5172 4632 5224 4684
rect 9588 4768 9640 4820
rect 11244 4768 11296 4820
rect 11520 4768 11572 4820
rect 5264 4607 5316 4616
rect 5264 4573 5273 4607
rect 5273 4573 5307 4607
rect 5307 4573 5316 4607
rect 5264 4564 5316 4573
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 7840 4564 7892 4616
rect 10968 4564 11020 4616
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 11612 4632 11664 4684
rect 11980 4632 12032 4684
rect 6368 4496 6420 4548
rect 7196 4496 7248 4548
rect 11704 4539 11756 4548
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 11704 4505 11713 4539
rect 11713 4505 11747 4539
rect 11747 4505 11756 4539
rect 12348 4607 12400 4616
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 13452 4768 13504 4820
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 14556 4768 14608 4820
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 12900 4564 12952 4616
rect 11704 4496 11756 4505
rect 13912 4428 13964 4480
rect 14648 4496 14700 4548
rect 14280 4471 14332 4480
rect 14280 4437 14307 4471
rect 14307 4437 14332 4471
rect 14280 4428 14332 4437
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 15200 4428 15252 4480
rect 15568 4428 15620 4480
rect 7214 4326 7266 4378
rect 7278 4326 7330 4378
rect 7342 4326 7394 4378
rect 7406 4326 7458 4378
rect 7470 4326 7522 4378
rect 13214 4326 13266 4378
rect 13278 4326 13330 4378
rect 13342 4326 13394 4378
rect 13406 4326 13458 4378
rect 13470 4326 13522 4378
rect 5816 4267 5868 4276
rect 5816 4233 5825 4267
rect 5825 4233 5859 4267
rect 5859 4233 5868 4267
rect 5816 4224 5868 4233
rect 6736 4224 6788 4276
rect 7104 4224 7156 4276
rect 7564 4224 7616 4276
rect 20 4088 72 4140
rect 3424 4156 3476 4208
rect 3516 4156 3568 4208
rect 5172 4156 5224 4208
rect 5632 4199 5684 4208
rect 5632 4165 5641 4199
rect 5641 4165 5675 4199
rect 5675 4165 5684 4199
rect 5632 4156 5684 4165
rect 6276 4156 6328 4208
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 8116 4199 8168 4208
rect 8116 4165 8125 4199
rect 8125 4165 8159 4199
rect 8159 4165 8168 4199
rect 8116 4156 8168 4165
rect 8484 4224 8536 4276
rect 11336 4224 11388 4276
rect 11520 4156 11572 4208
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 6460 3952 6512 4004
rect 8208 4020 8260 4072
rect 11152 4088 11204 4140
rect 11612 4088 11664 4140
rect 12348 4088 12400 4140
rect 13636 4224 13688 4276
rect 12716 4156 12768 4208
rect 13544 4156 13596 4208
rect 13912 4199 13964 4208
rect 13912 4165 13921 4199
rect 13921 4165 13955 4199
rect 13955 4165 13964 4199
rect 13912 4156 13964 4165
rect 14280 4156 14332 4208
rect 11428 4020 11480 4072
rect 11980 4020 12032 4072
rect 12992 4088 13044 4140
rect 8484 3952 8536 4004
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 12808 3927 12860 3936
rect 12808 3893 12817 3927
rect 12817 3893 12851 3927
rect 12851 3893 12860 3927
rect 12808 3884 12860 3893
rect 12992 3884 13044 3936
rect 13176 3884 13228 3936
rect 13912 3884 13964 3936
rect 15568 4156 15620 4208
rect 14740 4131 14792 4140
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 10214 3782 10266 3834
rect 10278 3782 10330 3834
rect 10342 3782 10394 3834
rect 10406 3782 10458 3834
rect 10470 3782 10522 3834
rect 16214 3782 16266 3834
rect 16278 3782 16330 3834
rect 16342 3782 16394 3834
rect 16406 3782 16458 3834
rect 16470 3782 16522 3834
rect 5172 3680 5224 3732
rect 6276 3723 6328 3732
rect 6276 3689 6285 3723
rect 6285 3689 6319 3723
rect 6319 3689 6328 3723
rect 6276 3680 6328 3689
rect 6368 3680 6420 3732
rect 6460 3680 6512 3732
rect 8484 3544 8536 3596
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 11152 3519 11204 3528
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 8116 3383 8168 3392
rect 8116 3349 8125 3383
rect 8125 3349 8159 3383
rect 8159 3349 8168 3383
rect 8116 3340 8168 3349
rect 10140 3340 10192 3392
rect 12072 3340 12124 3392
rect 12808 3680 12860 3732
rect 12900 3680 12952 3732
rect 14004 3680 14056 3732
rect 13084 3612 13136 3664
rect 12808 3544 12860 3596
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 12624 3451 12676 3460
rect 12624 3417 12633 3451
rect 12633 3417 12667 3451
rect 12667 3417 12676 3451
rect 12624 3408 12676 3417
rect 12992 3383 13044 3392
rect 12992 3349 13001 3383
rect 13001 3349 13035 3383
rect 13035 3349 13044 3383
rect 12992 3340 13044 3349
rect 13176 3383 13228 3392
rect 13176 3349 13203 3383
rect 13203 3349 13228 3383
rect 13176 3340 13228 3349
rect 13728 3476 13780 3528
rect 13912 3476 13964 3528
rect 13544 3408 13596 3460
rect 14280 3451 14332 3460
rect 14280 3417 14289 3451
rect 14289 3417 14323 3451
rect 14323 3417 14332 3451
rect 14280 3408 14332 3417
rect 15292 3340 15344 3392
rect 7214 3238 7266 3290
rect 7278 3238 7330 3290
rect 7342 3238 7394 3290
rect 7406 3238 7458 3290
rect 7470 3238 7522 3290
rect 13214 3238 13266 3290
rect 13278 3238 13330 3290
rect 13342 3238 13394 3290
rect 13406 3238 13458 3290
rect 13470 3238 13522 3290
rect 7104 3136 7156 3188
rect 8484 3136 8536 3188
rect 9588 3136 9640 3188
rect 7196 3000 7248 3052
rect 8484 3000 8536 3052
rect 10140 3068 10192 3120
rect 10968 3000 11020 3052
rect 11704 3136 11756 3188
rect 14740 3136 14792 3188
rect 12072 3068 12124 3120
rect 14280 3068 14332 3120
rect 15108 3068 15160 3120
rect 15292 3068 15344 3120
rect 13544 3000 13596 3052
rect 13636 3000 13688 3052
rect 12992 2932 13044 2984
rect 11152 2864 11204 2916
rect 8208 2796 8260 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 10214 2694 10266 2746
rect 10278 2694 10330 2746
rect 10342 2694 10394 2746
rect 10406 2694 10458 2746
rect 10470 2694 10522 2746
rect 16214 2694 16266 2746
rect 16278 2694 16330 2746
rect 16342 2694 16394 2746
rect 16406 2694 16458 2746
rect 16470 2694 16522 2746
rect 7196 2635 7248 2644
rect 7196 2601 7205 2635
rect 7205 2601 7239 2635
rect 7239 2601 7248 2635
rect 7196 2592 7248 2601
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 10600 2592 10652 2644
rect 11704 2635 11756 2644
rect 11704 2601 11713 2635
rect 11713 2601 11747 2635
rect 11747 2601 11756 2635
rect 11704 2592 11756 2601
rect 15384 2592 15436 2644
rect 7012 2388 7064 2440
rect 8116 2524 8168 2576
rect 8484 2567 8536 2576
rect 8484 2533 8493 2567
rect 8493 2533 8527 2567
rect 8527 2533 8536 2567
rect 8484 2524 8536 2533
rect 8392 2456 8444 2508
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 17040 2388 17092 2440
rect 4620 2363 4672 2372
rect 4620 2329 4629 2363
rect 4629 2329 4663 2363
rect 4663 2329 4672 2363
rect 4620 2320 4672 2329
rect 8208 2320 8260 2372
rect 7214 2150 7266 2202
rect 7278 2150 7330 2202
rect 7342 2150 7394 2202
rect 7406 2150 7458 2202
rect 7470 2150 7522 2202
rect 13214 2150 13266 2202
rect 13278 2150 13330 2202
rect 13342 2150 13394 2202
rect 13406 2150 13458 2202
rect 13470 2150 13522 2202
<< metal2 >>
rect 662 19650 718 20450
rect 5814 19650 5870 20450
rect 10966 19802 11022 20450
rect 10704 19774 11022 19802
rect 676 17746 704 19650
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 664 17740 716 17746
rect 664 17682 716 17688
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 1596 17202 1624 17478
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 1584 17196 1636 17202
rect 1584 17138 1636 17144
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2056 16574 2084 17138
rect 2608 16726 2636 17274
rect 2700 17134 2728 17478
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2884 16794 2912 17614
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2136 16584 2188 16590
rect 2056 16546 2136 16574
rect 2608 16574 2636 16662
rect 4080 16658 4108 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 2608 16546 2728 16574
rect 2136 16526 2188 16532
rect 2148 16114 2176 16526
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2240 16114 2268 16186
rect 2332 16114 2360 16458
rect 2700 16114 2728 16546
rect 5460 16522 5488 17138
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5552 16590 5580 16934
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5828 16538 5856 19650
rect 10214 17980 10522 17989
rect 10214 17978 10220 17980
rect 10276 17978 10300 17980
rect 10356 17978 10380 17980
rect 10436 17978 10460 17980
rect 10516 17978 10522 17980
rect 10276 17926 10278 17978
rect 10458 17926 10460 17978
rect 10214 17924 10220 17926
rect 10276 17924 10300 17926
rect 10356 17924 10380 17926
rect 10436 17924 10460 17926
rect 10516 17924 10522 17926
rect 10214 17915 10522 17924
rect 7214 17436 7522 17445
rect 7214 17434 7220 17436
rect 7276 17434 7300 17436
rect 7356 17434 7380 17436
rect 7436 17434 7460 17436
rect 7516 17434 7522 17436
rect 7276 17382 7278 17434
rect 7458 17382 7460 17434
rect 7214 17380 7220 17382
rect 7276 17380 7300 17382
rect 7356 17380 7380 17382
rect 7436 17380 7460 17382
rect 7516 17380 7522 17382
rect 7214 17371 7522 17380
rect 10704 17202 10732 19774
rect 10966 19650 11022 19774
rect 16118 19650 16174 20450
rect 16132 17762 16160 19650
rect 16214 17980 16522 17989
rect 16214 17978 16220 17980
rect 16276 17978 16300 17980
rect 16356 17978 16380 17980
rect 16436 17978 16460 17980
rect 16516 17978 16522 17980
rect 16276 17926 16278 17978
rect 16458 17926 16460 17978
rect 16214 17924 16220 17926
rect 16276 17924 16300 17926
rect 16356 17924 16380 17926
rect 16436 17924 16460 17926
rect 16516 17924 16522 17926
rect 16214 17915 16522 17924
rect 17038 17776 17094 17785
rect 16132 17734 16252 17762
rect 16224 17678 16252 17734
rect 17038 17711 17040 17720
rect 17092 17711 17094 17720
rect 17040 17682 17092 17688
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 13214 17436 13522 17445
rect 13214 17434 13220 17436
rect 13276 17434 13300 17436
rect 13356 17434 13380 17436
rect 13436 17434 13460 17436
rect 13516 17434 13522 17436
rect 13276 17382 13278 17434
rect 13458 17382 13460 17434
rect 13214 17380 13220 17382
rect 13276 17380 13300 17382
rect 13356 17380 13380 17382
rect 13436 17380 13460 17382
rect 13516 17380 13522 17382
rect 13214 17371 13522 17380
rect 15948 17338 15976 17478
rect 16224 17338 16252 17478
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11888 17128 11940 17134
rect 11888 17070 11940 17076
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 10214 16892 10522 16901
rect 10214 16890 10220 16892
rect 10276 16890 10300 16892
rect 10356 16890 10380 16892
rect 10436 16890 10460 16892
rect 10516 16890 10522 16892
rect 10276 16838 10278 16890
rect 10458 16838 10460 16890
rect 10214 16836 10220 16838
rect 10276 16836 10300 16838
rect 10356 16836 10380 16838
rect 10436 16836 10460 16838
rect 10516 16836 10522 16838
rect 10214 16827 10522 16836
rect 11256 16794 11284 16934
rect 11808 16794 11836 17070
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11428 16584 11480 16590
rect 5448 16516 5500 16522
rect 5828 16510 5948 16538
rect 11900 16574 11928 17070
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 11480 16546 11928 16574
rect 12544 16574 12572 16934
rect 12544 16546 12848 16574
rect 11428 16526 11480 16532
rect 5448 16458 5500 16464
rect 940 16108 992 16114
rect 940 16050 992 16056
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 952 15745 980 16050
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 938 15736 994 15745
rect 938 15671 994 15680
rect 1688 12306 1716 15846
rect 1780 15570 1808 15846
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 1780 15094 1808 15506
rect 1768 15088 1820 15094
rect 1768 15030 1820 15036
rect 2148 15026 2176 16050
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2240 14958 2268 16050
rect 2332 15026 2360 16050
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2700 15570 2728 15846
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2792 15026 2820 15914
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3344 15094 3372 15302
rect 3332 15088 3384 15094
rect 3332 15030 3384 15036
rect 4172 15026 4200 15370
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4816 15026 4844 15302
rect 5276 15026 5304 15846
rect 5460 15638 5488 16458
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5552 16250 5580 16390
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5828 16114 5856 16390
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5368 15162 5396 15438
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2516 12918 2544 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3988 14074 4016 14214
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3436 13326 3464 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 4632 13190 4660 14962
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14618 4844 14758
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 2504 12912 2556 12918
rect 2504 12854 2556 12860
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12434 3096 12582
rect 2884 12406 3096 12434
rect 3436 12434 3464 13126
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3436 12406 3556 12434
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 2136 12164 2188 12170
rect 2136 12106 2188 12112
rect 2148 11354 2176 12106
rect 2884 11762 2912 12406
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11898 3464 12038
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 940 10600 992 10606
rect 940 10542 992 10548
rect 952 10305 980 10542
rect 938 10296 994 10305
rect 938 10231 994 10240
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1872 9722 1900 9930
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1872 8974 1900 9522
rect 2424 9178 2452 11086
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2792 10146 2820 10610
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2872 10192 2924 10198
rect 2792 10140 2872 10146
rect 2792 10134 2924 10140
rect 2792 10118 2912 10134
rect 2792 9722 2820 10118
rect 3068 9722 3096 10202
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3160 9518 3188 9862
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 5370 1624 8774
rect 3344 8498 3372 10406
rect 3528 9602 3556 12406
rect 4632 12170 4660 13126
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 3712 9926 3740 12106
rect 4632 11830 4660 12106
rect 4724 11898 4752 12174
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4816 11762 4844 12582
rect 4908 11762 4936 12786
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5276 12238 5304 12650
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4080 11626 4200 11642
rect 4080 11620 4212 11626
rect 4080 11614 4160 11620
rect 4080 11150 4108 11614
rect 4160 11562 4212 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4080 10062 4108 11086
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4356 10810 4384 11018
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4632 10674 4660 11222
rect 4816 11150 4844 11698
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4724 10606 4752 10950
rect 4816 10810 4844 11086
rect 4908 11014 4936 11698
rect 5000 11150 5028 11698
rect 5736 11218 5764 12718
rect 5920 12714 5948 16510
rect 7214 16348 7522 16357
rect 7214 16346 7220 16348
rect 7276 16346 7300 16348
rect 7356 16346 7380 16348
rect 7436 16346 7460 16348
rect 7516 16346 7522 16348
rect 7276 16294 7278 16346
rect 7458 16294 7460 16346
rect 7214 16292 7220 16294
rect 7276 16292 7300 16294
rect 7356 16292 7380 16294
rect 7436 16292 7460 16294
rect 7516 16292 7522 16294
rect 7214 16283 7522 16292
rect 10214 15804 10522 15813
rect 10214 15802 10220 15804
rect 10276 15802 10300 15804
rect 10356 15802 10380 15804
rect 10436 15802 10460 15804
rect 10516 15802 10522 15804
rect 10276 15750 10278 15802
rect 10458 15750 10460 15802
rect 10214 15748 10220 15750
rect 10276 15748 10300 15750
rect 10356 15748 10380 15750
rect 10436 15748 10460 15750
rect 10516 15748 10522 15750
rect 10214 15739 10522 15748
rect 11440 15638 11468 16526
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12636 16114 12664 16390
rect 12728 16114 12756 16390
rect 12820 16114 12848 16546
rect 12912 16538 12940 17138
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 16794 13308 16934
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 12912 16522 13308 16538
rect 12912 16516 13320 16522
rect 12912 16510 13268 16516
rect 13268 16458 13320 16464
rect 13372 16454 13400 17070
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16590 13860 16934
rect 16214 16892 16522 16901
rect 16214 16890 16220 16892
rect 16276 16890 16300 16892
rect 16356 16890 16380 16892
rect 16436 16890 16460 16892
rect 16516 16890 16522 16892
rect 16276 16838 16278 16890
rect 16458 16838 16460 16890
rect 16214 16836 16220 16838
rect 16276 16836 16300 16838
rect 16356 16836 16380 16838
rect 16436 16836 16460 16838
rect 16516 16836 16522 16838
rect 16214 16827 16522 16836
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13214 16348 13522 16357
rect 13214 16346 13220 16348
rect 13276 16346 13300 16348
rect 13356 16346 13380 16348
rect 13436 16346 13460 16348
rect 13516 16346 13522 16348
rect 13276 16294 13278 16346
rect 13458 16294 13460 16346
rect 13214 16292 13220 16294
rect 13276 16292 13300 16294
rect 13356 16292 13380 16294
rect 13436 16292 13460 16294
rect 13516 16292 13522 16294
rect 13214 16283 13522 16292
rect 13556 16182 13584 16390
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 6104 15026 6132 15370
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7116 15094 7144 15302
rect 7214 15260 7522 15269
rect 7214 15258 7220 15260
rect 7276 15258 7300 15260
rect 7356 15258 7380 15260
rect 7436 15258 7460 15260
rect 7516 15258 7522 15260
rect 7276 15206 7278 15258
rect 7458 15206 7460 15258
rect 7214 15204 7220 15206
rect 7276 15204 7300 15206
rect 7356 15204 7380 15206
rect 7436 15204 7460 15206
rect 7516 15204 7522 15206
rect 7214 15195 7522 15204
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 8312 15026 8340 15370
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8496 15094 8524 15302
rect 8680 15162 8708 15370
rect 9048 15162 9076 15438
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 8484 15088 8536 15094
rect 8484 15030 8536 15036
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 6840 14618 6868 14962
rect 8496 14618 8524 15030
rect 8680 15026 8708 15098
rect 9048 15026 9076 15098
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8956 14414 8984 14962
rect 9324 14482 9352 15302
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7214 14172 7522 14181
rect 7214 14170 7220 14172
rect 7276 14170 7300 14172
rect 7356 14170 7380 14172
rect 7436 14170 7460 14172
rect 7516 14170 7522 14172
rect 7276 14118 7278 14170
rect 7458 14118 7460 14170
rect 7214 14116 7220 14118
rect 7276 14116 7300 14118
rect 7356 14116 7380 14118
rect 7436 14116 7460 14118
rect 7516 14116 7522 14118
rect 7214 14107 7522 14116
rect 7852 14074 7880 14282
rect 8956 14074 8984 14350
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9416 14006 9444 14758
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9416 13394 9444 13942
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6288 12850 6316 13262
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 3712 9654 3740 9862
rect 3436 9574 3556 9602
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 4448 9602 4476 9862
rect 4540 9722 4568 9862
rect 4632 9722 4660 10134
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4724 9602 4752 10542
rect 4816 10062 4844 10746
rect 5000 10062 5028 11086
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5552 10266 5580 10610
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5828 10062 5856 10950
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5920 9738 5948 12650
rect 6288 12374 6316 12786
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6472 12238 6500 12582
rect 6564 12442 6592 13194
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7214 13084 7522 13093
rect 7214 13082 7220 13084
rect 7276 13082 7300 13084
rect 7356 13082 7380 13084
rect 7436 13082 7460 13084
rect 7516 13082 7522 13084
rect 7276 13030 7278 13082
rect 7458 13030 7460 13082
rect 7214 13028 7220 13030
rect 7276 13028 7300 13030
rect 7356 13028 7380 13030
rect 7436 13028 7460 13030
rect 7516 13028 7522 13030
rect 7214 13019 7522 13028
rect 8036 12986 8064 13126
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8312 12918 8340 13194
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6656 11762 6684 12650
rect 6932 11898 6960 12718
rect 7116 12374 7144 12786
rect 7104 12368 7156 12374
rect 7104 12310 7156 12316
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7116 11830 7144 12310
rect 7214 11996 7522 12005
rect 7214 11994 7220 11996
rect 7276 11994 7300 11996
rect 7356 11994 7380 11996
rect 7436 11994 7460 11996
rect 7516 11994 7522 11996
rect 7276 11942 7278 11994
rect 7458 11942 7460 11994
rect 7214 11940 7220 11942
rect 7276 11940 7300 11942
rect 7356 11940 7380 11942
rect 7436 11940 7460 11942
rect 7516 11940 7522 11942
rect 7214 11931 7522 11940
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7024 11354 7052 11494
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6012 10810 6040 11086
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6288 10674 6316 10950
rect 6840 10742 6868 11086
rect 7214 10908 7522 10917
rect 7214 10906 7220 10908
rect 7276 10906 7300 10908
rect 7356 10906 7380 10908
rect 7436 10906 7460 10908
rect 7516 10906 7522 10908
rect 7276 10854 7278 10906
rect 7458 10854 7460 10906
rect 7214 10852 7220 10854
rect 7276 10852 7300 10854
rect 7356 10852 7380 10854
rect 7436 10852 7460 10854
rect 7516 10852 7522 10854
rect 7214 10843 7522 10852
rect 7668 10810 7696 11698
rect 8864 11558 8892 13194
rect 9324 12986 9352 13194
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9416 12866 9444 13330
rect 9416 12850 9536 12866
rect 9416 12844 9548 12850
rect 9416 12838 9496 12844
rect 9496 12786 9548 12792
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 11762 9168 12582
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 7944 11354 7972 11494
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 8864 11082 8892 11494
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 8680 10742 8708 10950
rect 8864 10742 8892 11018
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6288 10062 6316 10610
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6288 9926 6316 9998
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 4448 9574 4752 9602
rect 5828 9710 5948 9738
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3436 7886 3464 9574
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7546 2820 7686
rect 4632 7546 4660 9574
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8906 4936 9318
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5000 8634 5028 8842
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5828 8498 5856 9710
rect 6288 9110 6316 9862
rect 6380 9674 6408 9998
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7214 9820 7522 9829
rect 7214 9818 7220 9820
rect 7276 9818 7300 9820
rect 7356 9818 7380 9820
rect 7436 9818 7460 9820
rect 7516 9818 7522 9820
rect 7276 9766 7278 9818
rect 7458 9766 7460 9818
rect 7214 9764 7220 9766
rect 7276 9764 7300 9766
rect 7356 9764 7380 9766
rect 7436 9764 7460 9766
rect 7516 9764 7522 9766
rect 7214 9755 7522 9764
rect 6380 9646 6500 9674
rect 6472 9382 6500 9646
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6104 8566 6132 8910
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5828 8362 5856 8434
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 6104 7750 6132 8502
rect 6288 7954 6316 9046
rect 6472 9042 6500 9318
rect 7668 9110 7696 9318
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7760 9042 7788 9862
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 6472 8566 6500 8774
rect 7214 8732 7522 8741
rect 7214 8730 7220 8732
rect 7276 8730 7300 8732
rect 7356 8730 7380 8732
rect 7436 8730 7460 8732
rect 7516 8730 7522 8732
rect 7276 8678 7278 8730
rect 7458 8678 7460 8730
rect 7214 8676 7220 8678
rect 7276 8676 7300 8678
rect 7356 8676 7380 8678
rect 7436 8676 7460 8678
rect 7516 8676 7522 8678
rect 7214 8667 7522 8676
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 7576 8430 7604 8774
rect 7760 8634 7788 8774
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 8588 8566 8616 9590
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 9178 9536 9454
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7954 6960 8230
rect 8404 8090 8432 8502
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 8588 7818 8616 8502
rect 9600 7886 9628 14962
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9692 11830 9720 14826
rect 10214 14716 10522 14725
rect 10214 14714 10220 14716
rect 10276 14714 10300 14716
rect 10356 14714 10380 14716
rect 10436 14714 10460 14716
rect 10516 14714 10522 14716
rect 10276 14662 10278 14714
rect 10458 14662 10460 14714
rect 10214 14660 10220 14662
rect 10276 14660 10300 14662
rect 10356 14660 10380 14662
rect 10436 14660 10460 14662
rect 10516 14660 10522 14662
rect 10214 14651 10522 14660
rect 10704 14346 10732 15098
rect 10980 15094 11008 15370
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10980 14414 11008 15030
rect 11348 14958 11376 15302
rect 11440 15026 11468 15302
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11072 14618 11100 14894
rect 11440 14618 11468 14962
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11624 14482 11652 14962
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 12268 14414 12296 14554
rect 12452 14550 12480 14758
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9876 12646 9904 12786
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 10152 12306 10180 13806
rect 10214 13628 10522 13637
rect 10214 13626 10220 13628
rect 10276 13626 10300 13628
rect 10356 13626 10380 13628
rect 10436 13626 10460 13628
rect 10516 13626 10522 13628
rect 10276 13574 10278 13626
rect 10458 13574 10460 13626
rect 10214 13572 10220 13574
rect 10276 13572 10300 13574
rect 10356 13572 10380 13574
rect 10436 13572 10460 13574
rect 10516 13572 10522 13574
rect 10214 13563 10522 13572
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10428 12850 10456 13330
rect 10704 13326 10732 14282
rect 12268 13870 12296 14350
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10612 12714 10640 12922
rect 10796 12850 10824 12922
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10214 12540 10522 12549
rect 10214 12538 10220 12540
rect 10276 12538 10300 12540
rect 10356 12538 10380 12540
rect 10436 12538 10460 12540
rect 10516 12538 10522 12540
rect 10276 12486 10278 12538
rect 10458 12486 10460 12538
rect 10214 12484 10220 12486
rect 10276 12484 10300 12486
rect 10356 12484 10380 12486
rect 10436 12484 10460 12486
rect 10516 12484 10522 12486
rect 10214 12475 10522 12484
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9876 10810 9904 11698
rect 10214 11452 10522 11461
rect 10214 11450 10220 11452
rect 10276 11450 10300 11452
rect 10356 11450 10380 11452
rect 10436 11450 10460 11452
rect 10516 11450 10522 11452
rect 10276 11398 10278 11450
rect 10458 11398 10460 11450
rect 10214 11396 10220 11398
rect 10276 11396 10300 11398
rect 10356 11396 10380 11398
rect 10436 11396 10460 11398
rect 10516 11396 10522 11398
rect 10214 11387 10522 11396
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10152 10810 10180 11018
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10214 10364 10522 10373
rect 10214 10362 10220 10364
rect 10276 10362 10300 10364
rect 10356 10362 10380 10364
rect 10436 10362 10460 10364
rect 10516 10362 10522 10364
rect 10276 10310 10278 10362
rect 10458 10310 10460 10362
rect 10214 10308 10220 10310
rect 10276 10308 10300 10310
rect 10356 10308 10380 10310
rect 10436 10308 10460 10310
rect 10516 10308 10522 10310
rect 10214 10299 10522 10308
rect 10214 9276 10522 9285
rect 10214 9274 10220 9276
rect 10276 9274 10300 9276
rect 10356 9274 10380 9276
rect 10436 9274 10460 9276
rect 10516 9274 10522 9276
rect 10276 9222 10278 9274
rect 10458 9222 10460 9274
rect 10214 9220 10220 9222
rect 10276 9220 10300 9222
rect 10356 9220 10380 9222
rect 10436 9220 10460 9222
rect 10516 9220 10522 9222
rect 10214 9211 10522 9220
rect 10214 8188 10522 8197
rect 10214 8186 10220 8188
rect 10276 8186 10300 8188
rect 10356 8186 10380 8188
rect 10436 8186 10460 8188
rect 10516 8186 10522 8188
rect 10276 8134 10278 8186
rect 10458 8134 10460 8186
rect 10214 8132 10220 8134
rect 10276 8132 10300 8134
rect 10356 8132 10380 8134
rect 10436 8132 10460 8134
rect 10516 8132 10522 8134
rect 10214 8123 10522 8132
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 6104 7478 6132 7686
rect 7214 7644 7522 7653
rect 7214 7642 7220 7644
rect 7276 7642 7300 7644
rect 7356 7642 7380 7644
rect 7436 7642 7460 7644
rect 7516 7642 7522 7644
rect 7276 7590 7278 7642
rect 7458 7590 7460 7642
rect 7214 7588 7220 7590
rect 7276 7588 7300 7590
rect 7356 7588 7380 7590
rect 7436 7588 7460 7590
rect 7516 7588 7522 7590
rect 7214 7579 7522 7588
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 3620 6322 3648 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6322 4660 7142
rect 6012 7002 6040 7142
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2700 5914 2728 6190
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 5000 5914 5028 6258
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4865 980 5170
rect 938 4856 994 4865
rect 938 4791 994 4800
rect 3436 4214 3464 5578
rect 4908 5370 4936 5646
rect 5184 5574 5212 6326
rect 7024 6322 7052 6598
rect 7214 6556 7522 6565
rect 7214 6554 7220 6556
rect 7276 6554 7300 6556
rect 7356 6554 7380 6556
rect 7436 6554 7460 6556
rect 7516 6554 7522 6556
rect 7276 6502 7278 6554
rect 7458 6502 7460 6554
rect 7214 6500 7220 6502
rect 7276 6500 7300 6502
rect 7356 6500 7380 6502
rect 7436 6500 7460 6502
rect 7516 6500 7522 6502
rect 7214 6491 7522 6500
rect 7668 6322 7696 6802
rect 8128 6662 8156 6802
rect 8220 6730 8248 7686
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5828 5778 5856 6054
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3528 4214 3556 5102
rect 4080 4826 4108 5170
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 5184 4690 5212 5510
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5356 5228 5408 5234
rect 5408 5188 5580 5216
rect 5356 5170 5408 5176
rect 5552 5030 5580 5188
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 4214 5212 4626
rect 5276 4622 5304 4966
rect 5644 4826 5672 5238
rect 5828 5030 5856 5714
rect 7852 5574 7880 6326
rect 8036 5710 8064 6598
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7214 5468 7522 5477
rect 7214 5466 7220 5468
rect 7276 5466 7300 5468
rect 7356 5466 7380 5468
rect 7436 5466 7460 5468
rect 7516 5466 7522 5468
rect 7276 5414 7278 5466
rect 7458 5414 7460 5466
rect 7214 5412 7220 5414
rect 7276 5412 7300 5414
rect 7356 5412 7380 5414
rect 7436 5412 7460 5414
rect 7516 5412 7522 5414
rect 7214 5403 7522 5412
rect 7852 5234 7880 5510
rect 8036 5302 8064 5646
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5644 4214 5672 4762
rect 5828 4282 5856 4966
rect 6380 4554 6408 4966
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 20 4140 72 4146
rect 20 4082 72 4088
rect 32 800 60 4082
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5184 3738 5212 4150
rect 6288 3738 6316 4150
rect 6380 4146 6408 4490
rect 6748 4486 6776 4966
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6748 4282 6776 4422
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3738 6408 3878
rect 6472 3738 6500 3946
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7024 2446 7052 4762
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7116 4282 7144 4558
rect 7208 4554 7236 4966
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7214 4380 7522 4389
rect 7214 4378 7220 4380
rect 7276 4378 7300 4380
rect 7356 4378 7380 4380
rect 7436 4378 7460 4380
rect 7516 4378 7522 4380
rect 7276 4326 7278 4378
rect 7458 4326 7460 4378
rect 7214 4324 7220 4326
rect 7276 4324 7300 4326
rect 7356 4324 7380 4326
rect 7436 4324 7460 4326
rect 7516 4324 7522 4326
rect 7214 4315 7522 4324
rect 7576 4282 7604 5034
rect 7852 4622 7880 5170
rect 8128 5166 8156 6598
rect 8220 5166 8248 6666
rect 8772 6458 8800 6734
rect 9508 6662 9536 7346
rect 9600 7002 9628 7822
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7546 9812 7754
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 9508 6254 9536 6598
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9600 5574 9628 6938
rect 9692 6934 9720 7346
rect 10214 7100 10522 7109
rect 10214 7098 10220 7100
rect 10276 7098 10300 7100
rect 10356 7098 10380 7100
rect 10436 7098 10460 7100
rect 10516 7098 10522 7100
rect 10276 7046 10278 7098
rect 10458 7046 10460 7098
rect 10214 7044 10220 7046
rect 10276 7044 10300 7046
rect 10356 7044 10380 7046
rect 10436 7044 10460 7046
rect 10516 7044 10522 7046
rect 10214 7035 10522 7044
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 5710 9996 6598
rect 10152 6458 10180 6802
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 6458 10456 6666
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10214 6012 10522 6021
rect 10214 6010 10220 6012
rect 10276 6010 10300 6012
rect 10356 6010 10380 6012
rect 10436 6010 10460 6012
rect 10516 6010 10522 6012
rect 10276 5958 10278 6010
rect 10458 5958 10460 6010
rect 10214 5956 10220 5958
rect 10276 5956 10300 5958
rect 10356 5956 10380 5958
rect 10436 5956 10460 5958
rect 10516 5956 10522 5958
rect 10214 5947 10522 5956
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7116 3194 7144 4218
rect 8128 4214 8156 5102
rect 8220 4826 8248 5102
rect 9600 4826 9628 5510
rect 9784 5166 9812 5646
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 10214 4924 10522 4933
rect 10214 4922 10220 4924
rect 10276 4922 10300 4924
rect 10356 4922 10380 4924
rect 10436 4922 10460 4924
rect 10516 4922 10522 4924
rect 10276 4870 10278 4922
rect 10458 4870 10460 4922
rect 10214 4868 10220 4870
rect 10276 4868 10300 4870
rect 10356 4868 10380 4870
rect 10436 4868 10460 4870
rect 10516 4868 10522 4870
rect 10214 4859 10522 4868
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8496 4282 8524 4422
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7214 3292 7522 3301
rect 7214 3290 7220 3292
rect 7276 3290 7300 3292
rect 7356 3290 7380 3292
rect 7436 3290 7460 3292
rect 7516 3290 7522 3292
rect 7276 3238 7278 3290
rect 7458 3238 7460 3290
rect 7214 3236 7220 3238
rect 7276 3236 7300 3238
rect 7356 3236 7380 3238
rect 7436 3236 7460 3238
rect 7516 3236 7522 3238
rect 7214 3227 7522 3236
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7208 2650 7236 2994
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 8128 2582 8156 3334
rect 8220 2854 8248 4014
rect 8496 4010 8524 4082
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8496 3602 8524 3946
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 8220 2378 8248 2790
rect 8404 2514 8432 3470
rect 8496 3194 8524 3538
rect 9600 3194 9628 4762
rect 10214 3836 10522 3845
rect 10214 3834 10220 3836
rect 10276 3834 10300 3836
rect 10356 3834 10380 3836
rect 10436 3834 10460 3836
rect 10516 3834 10522 3836
rect 10276 3782 10278 3834
rect 10458 3782 10460 3834
rect 10214 3780 10220 3782
rect 10276 3780 10300 3782
rect 10356 3780 10380 3782
rect 10436 3780 10460 3782
rect 10516 3780 10522 3782
rect 10214 3771 10522 3780
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8496 2582 8524 2994
rect 9600 2774 9628 3130
rect 10152 3126 10180 3334
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 9508 2746 9628 2774
rect 10214 2748 10522 2757
rect 10214 2746 10220 2748
rect 10276 2746 10300 2748
rect 10356 2746 10380 2748
rect 10436 2746 10460 2748
rect 10516 2746 10522 2748
rect 9508 2650 9536 2746
rect 10276 2694 10278 2746
rect 10458 2694 10460 2746
rect 10214 2692 10220 2694
rect 10276 2692 10300 2694
rect 10356 2692 10380 2694
rect 10436 2692 10460 2694
rect 10516 2692 10522 2694
rect 10214 2683 10522 2692
rect 10612 2650 10640 12650
rect 10888 12434 10916 13126
rect 12452 12918 12480 13262
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12268 12442 12296 12582
rect 10796 12406 10916 12434
rect 12256 12436 12308 12442
rect 10796 12306 10824 12406
rect 12256 12378 12308 12384
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 12452 12170 12480 12854
rect 12544 12782 12572 15846
rect 12820 14822 12848 16050
rect 13096 15706 13124 16050
rect 14200 16046 14228 16526
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13214 15260 13522 15269
rect 13214 15258 13220 15260
rect 13276 15258 13300 15260
rect 13356 15258 13380 15260
rect 13436 15258 13460 15260
rect 13516 15258 13522 15260
rect 13276 15206 13278 15258
rect 13458 15206 13460 15258
rect 13214 15204 13220 15206
rect 13276 15204 13300 15206
rect 13356 15204 13380 15206
rect 13436 15204 13460 15206
rect 13516 15204 13522 15206
rect 13214 15195 13522 15204
rect 14200 15162 14228 15982
rect 14292 15706 14320 16390
rect 14568 16114 14596 16458
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14568 15434 14596 16050
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15570 15516 15846
rect 16214 15804 16522 15813
rect 16214 15802 16220 15804
rect 16276 15802 16300 15804
rect 16356 15802 16380 15804
rect 16436 15802 16460 15804
rect 16516 15802 16522 15804
rect 16276 15750 16278 15802
rect 16458 15750 16460 15802
rect 16214 15748 16220 15750
rect 16276 15748 16300 15750
rect 16356 15748 16380 15750
rect 16436 15748 16460 15750
rect 16516 15748 16522 15750
rect 16214 15739 16522 15748
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13004 13938 13032 14758
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 14074 13124 14282
rect 13214 14172 13522 14181
rect 13214 14170 13220 14172
rect 13276 14170 13300 14172
rect 13356 14170 13380 14172
rect 13436 14170 13460 14172
rect 13516 14170 13522 14172
rect 13276 14118 13278 14170
rect 13458 14118 13460 14170
rect 13214 14116 13220 14118
rect 13276 14116 13300 14118
rect 13356 14116 13380 14118
rect 13436 14116 13460 14118
rect 13516 14116 13522 14118
rect 13214 14107 13522 14116
rect 13556 14074 13584 14758
rect 13832 14618 13860 15030
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13004 13410 13032 13874
rect 14292 13734 14320 14214
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 13004 13382 13124 13410
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12544 12374 12572 12718
rect 13096 12374 13124 13382
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13214 13084 13522 13093
rect 13214 13082 13220 13084
rect 13276 13082 13300 13084
rect 13356 13082 13380 13084
rect 13436 13082 13460 13084
rect 13516 13082 13522 13084
rect 13276 13030 13278 13082
rect 13458 13030 13460 13082
rect 13214 13028 13220 13030
rect 13276 13028 13300 13030
rect 13356 13028 13380 13030
rect 13436 13028 13460 13030
rect 13516 13028 13522 13030
rect 13214 13019 13522 13028
rect 13556 12986 13584 13194
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13832 12442 13860 13262
rect 14292 12646 14320 13670
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11164 11354 11192 11562
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11348 11354 11376 11494
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11164 10062 11192 11290
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11256 10198 11284 10542
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10888 8650 10916 9522
rect 10980 8974 11008 9930
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9382 11192 9862
rect 11256 9722 11284 10134
rect 11348 9722 11376 10134
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11440 9178 11468 11494
rect 12452 11218 12480 12106
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 11762 12756 12038
rect 13096 11898 13124 12310
rect 14292 12238 14320 12582
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13214 11996 13522 12005
rect 13214 11994 13220 11996
rect 13276 11994 13300 11996
rect 13356 11994 13380 11996
rect 13436 11994 13460 11996
rect 13516 11994 13522 11996
rect 13276 11942 13278 11994
rect 13458 11942 13460 11994
rect 13214 11940 13220 11942
rect 13276 11940 13300 11942
rect 13356 11940 13380 11942
rect 13436 11940 13460 11942
rect 13516 11940 13522 11942
rect 13214 11931 13522 11940
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12452 11082 12480 11154
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 10062 11560 10406
rect 12268 10130 12296 10678
rect 12636 10266 12664 10950
rect 12820 10656 12848 11698
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11354 13308 11494
rect 13556 11354 13584 11698
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13740 11150 13768 12106
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11898 14228 12038
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14292 11830 14320 12174
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 12900 10668 12952 10674
rect 12820 10628 12900 10656
rect 12900 10610 12952 10616
rect 12912 10266 12940 10610
rect 13096 10606 13124 11086
rect 13214 10908 13522 10917
rect 13214 10906 13220 10908
rect 13276 10906 13300 10908
rect 13356 10906 13380 10908
rect 13436 10906 13460 10908
rect 13516 10906 13522 10908
rect 13276 10854 13278 10906
rect 13458 10854 13460 10906
rect 13214 10852 13220 10854
rect 13276 10852 13300 10854
rect 13356 10852 13380 10854
rect 13436 10852 13460 10854
rect 13516 10852 13522 10854
rect 13214 10843 13522 10852
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 12268 9722 12296 10066
rect 13372 10062 13400 10406
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 12544 9722 12572 9930
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13214 9820 13522 9829
rect 13214 9818 13220 9820
rect 13276 9818 13300 9820
rect 13356 9818 13380 9820
rect 13436 9818 13460 9820
rect 13516 9818 13522 9820
rect 13276 9766 13278 9818
rect 13458 9766 13460 9818
rect 13214 9764 13220 9766
rect 13276 9764 13300 9766
rect 13356 9764 13380 9766
rect 13436 9764 13460 9766
rect 13516 9764 13522 9766
rect 13214 9755 13522 9764
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 13648 9602 13676 9862
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13556 9574 13676 9602
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10888 8622 11008 8650
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10888 8090 10916 8434
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10888 6882 10916 8026
rect 10980 7478 11008 8622
rect 11440 8498 11468 9114
rect 13096 8906 13124 9522
rect 13556 9518 13584 9574
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13924 9178 13952 9930
rect 14016 9654 14044 10542
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 9722 14228 10406
rect 14384 10266 14412 15370
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 14648 13932 14700 13938
rect 14648 13874 14700 13880
rect 14660 13530 14688 13874
rect 15304 13530 15332 14894
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14414 15608 14758
rect 15948 14618 15976 14962
rect 16214 14716 16522 14725
rect 16214 14714 16220 14716
rect 16276 14714 16300 14716
rect 16356 14714 16380 14716
rect 16436 14714 16460 14716
rect 16516 14714 16522 14716
rect 16276 14662 16278 14714
rect 16458 14662 16460 14714
rect 16214 14660 16220 14662
rect 16276 14660 16300 14662
rect 16356 14660 16380 14662
rect 16436 14660 16460 14662
rect 16516 14660 16522 14662
rect 16214 14651 16522 14660
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15488 13326 15516 14010
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15580 13326 15608 13670
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15568 13320 15620 13326
rect 15568 13262 15620 13268
rect 16040 13190 16068 13874
rect 16214 13628 16522 13637
rect 16214 13626 16220 13628
rect 16276 13626 16300 13628
rect 16356 13626 16380 13628
rect 16436 13626 16460 13628
rect 16516 13626 16522 13628
rect 16276 13574 16278 13626
rect 16458 13574 16460 13626
rect 16214 13572 16220 13574
rect 16276 13572 16300 13574
rect 16356 13572 16380 13574
rect 16436 13572 16460 13574
rect 16516 13572 16522 13574
rect 16214 13563 16522 13572
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15028 12322 15056 12854
rect 14936 12306 15056 12322
rect 14924 12300 15056 12306
rect 14976 12294 15056 12300
rect 14924 12242 14976 12248
rect 15028 11558 15056 12294
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15028 11082 15056 11494
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15120 10826 15148 11834
rect 15212 11218 15240 12854
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15304 12170 15332 12582
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15304 11354 15332 11698
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15120 10798 15240 10826
rect 15212 10674 15240 10798
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 14476 9382 14504 9862
rect 14752 9602 14780 9998
rect 14844 9722 14872 10610
rect 15120 9926 15148 10610
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14752 9574 14872 9602
rect 15488 9586 15516 10610
rect 15856 10606 15884 12786
rect 16040 12646 16068 13126
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16040 12220 16068 12582
rect 16132 12345 16160 12582
rect 16214 12540 16522 12549
rect 16214 12538 16220 12540
rect 16276 12538 16300 12540
rect 16356 12538 16380 12540
rect 16436 12538 16460 12540
rect 16516 12538 16522 12540
rect 16276 12486 16278 12538
rect 16458 12486 16460 12538
rect 16214 12484 16220 12486
rect 16276 12484 16300 12486
rect 16356 12484 16380 12486
rect 16436 12484 16460 12486
rect 16516 12484 16522 12486
rect 16214 12475 16522 12484
rect 16118 12336 16174 12345
rect 16118 12271 16174 12280
rect 16212 12232 16264 12238
rect 16040 12192 16212 12220
rect 16212 12174 16264 12180
rect 16214 11452 16522 11461
rect 16214 11450 16220 11452
rect 16276 11450 16300 11452
rect 16356 11450 16380 11452
rect 16436 11450 16460 11452
rect 16516 11450 16522 11452
rect 16276 11398 16278 11450
rect 16458 11398 16460 11450
rect 16214 11396 16220 11398
rect 16276 11396 16300 11398
rect 16356 11396 16380 11398
rect 16436 11396 16460 11398
rect 16516 11396 16522 11398
rect 16214 11387 16522 11396
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 16214 10364 16522 10373
rect 16214 10362 16220 10364
rect 16276 10362 16300 10364
rect 16356 10362 16380 10364
rect 16436 10362 16460 10364
rect 16516 10362 16522 10364
rect 16276 10310 16278 10362
rect 16458 10310 16460 10362
rect 16214 10308 16220 10310
rect 16276 10308 16300 10310
rect 16356 10308 16380 10310
rect 16436 10308 16460 10310
rect 16516 10308 16522 10310
rect 16214 10299 16522 10308
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8634 13124 8842
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13214 8732 13522 8741
rect 13214 8730 13220 8732
rect 13276 8730 13300 8732
rect 13356 8730 13380 8732
rect 13436 8730 13460 8732
rect 13516 8730 13522 8732
rect 13276 8678 13278 8730
rect 13458 8678 13460 8730
rect 13214 8676 13220 8678
rect 13276 8676 13300 8678
rect 13356 8676 13380 8678
rect 13436 8676 13460 8678
rect 13516 8676 13522 8678
rect 13214 8667 13522 8676
rect 13556 8634 13584 8774
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11256 7886 11284 8298
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11440 7546 11468 8434
rect 11624 8090 11652 8434
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 13372 7834 13400 8298
rect 13648 8090 13676 8978
rect 13924 8498 13952 9114
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14384 8634 14412 8910
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13372 7806 13584 7834
rect 13214 7644 13522 7653
rect 13214 7642 13220 7644
rect 13276 7642 13300 7644
rect 13356 7642 13380 7644
rect 13436 7642 13460 7644
rect 13516 7642 13522 7644
rect 13276 7590 13278 7642
rect 13458 7590 13460 7642
rect 13214 7588 13220 7590
rect 13276 7588 13300 7590
rect 13356 7588 13380 7590
rect 13436 7588 13460 7590
rect 13516 7588 13522 7590
rect 13214 7579 13522 7588
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10796 6854 10916 6882
rect 10796 6662 10824 6854
rect 10980 6730 11008 7414
rect 11440 7410 11468 7482
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11440 6934 11468 7346
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 5642 10824 6598
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10980 4622 11008 6666
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11164 5914 11192 6258
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11900 5778 11928 6598
rect 11992 6458 12020 6598
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 12084 5710 12112 6802
rect 12268 6458 12296 7278
rect 12728 7002 12756 7414
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12360 6662 12388 6802
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12256 6248 12308 6254
rect 12452 6236 12480 6802
rect 12912 6322 12940 6870
rect 13004 6730 13032 7142
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 12900 6316 12952 6322
rect 12900 6258 12952 6264
rect 12308 6208 12480 6236
rect 12256 6190 12308 6196
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11072 5370 11100 5510
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11624 5302 11652 5510
rect 12084 5302 12112 5646
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11256 4826 11284 5102
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11532 4826 11560 5034
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 10980 3058 11008 4558
rect 11348 4282 11376 4558
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11532 4214 11560 4762
rect 11624 4690 11652 5238
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11716 4554 11744 5170
rect 11992 4690 12020 5170
rect 12176 5030 12204 6122
rect 12268 5710 12296 6190
rect 13004 6186 13032 6666
rect 13214 6556 13522 6565
rect 13214 6554 13220 6556
rect 13276 6554 13300 6556
rect 13356 6554 13380 6556
rect 13436 6554 13460 6556
rect 13516 6554 13522 6556
rect 13276 6502 13278 6554
rect 13458 6502 13460 6554
rect 13214 6500 13220 6502
rect 13276 6500 13300 6502
rect 13356 6500 13380 6502
rect 13436 6500 13460 6502
rect 13516 6500 13522 6502
rect 13214 6491 13522 6500
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12268 5302 12296 5646
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11704 4548 11756 4554
rect 11704 4490 11756 4496
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11164 3534 11192 4082
rect 11428 4072 11480 4078
rect 11624 4026 11652 4082
rect 11992 4078 12020 4626
rect 12360 4622 12388 5578
rect 12544 4622 12572 5714
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12820 5302 12848 5646
rect 13214 5468 13522 5477
rect 13214 5466 13220 5468
rect 13276 5466 13300 5468
rect 13356 5466 13380 5468
rect 13436 5466 13460 5468
rect 13516 5466 13522 5468
rect 13276 5414 13278 5466
rect 13458 5414 13460 5466
rect 13214 5412 13220 5414
rect 13276 5412 13300 5414
rect 13356 5412 13380 5414
rect 13436 5412 13460 5414
rect 13516 5412 13522 5414
rect 13214 5403 13522 5412
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12360 4146 12388 4558
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 11428 4014 11480 4020
rect 11440 3534 11468 4014
rect 11532 3998 11652 4026
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11532 3534 11560 3998
rect 12728 3618 12756 4150
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12820 3738 12848 3878
rect 12912 3738 12940 4558
rect 13004 4146 13032 4966
rect 13280 4690 13308 4966
rect 13556 4826 13584 7806
rect 13740 7546 13768 8434
rect 13832 7886 13860 8434
rect 14384 7954 14412 8570
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13648 6474 13676 6938
rect 13740 6798 13768 7482
rect 14568 7478 14596 8230
rect 14752 8090 14780 8230
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13648 6458 13952 6474
rect 13648 6452 13964 6458
rect 13648 6446 13912 6452
rect 13912 6394 13964 6400
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13648 5914 13676 6258
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13924 5642 13952 6054
rect 14752 5778 14780 6054
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14752 5658 14780 5714
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 14660 5630 14780 5658
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13832 5234 13860 5510
rect 14660 5302 14688 5630
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13464 4468 13492 4762
rect 13464 4440 13584 4468
rect 13214 4380 13522 4389
rect 13214 4378 13220 4380
rect 13276 4378 13300 4380
rect 13356 4378 13380 4380
rect 13436 4378 13460 4380
rect 13516 4378 13522 4380
rect 13276 4326 13278 4378
rect 13458 4326 13460 4378
rect 13214 4324 13220 4326
rect 13276 4324 13300 4326
rect 13356 4324 13380 4326
rect 13436 4324 13460 4326
rect 13516 4324 13522 4326
rect 13214 4315 13522 4324
rect 13556 4214 13584 4440
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12636 3590 12756 3618
rect 12820 3602 12848 3674
rect 12808 3596 12860 3602
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11164 2922 11192 3470
rect 12636 3466 12664 3590
rect 12808 3538 12860 3544
rect 12912 3534 12940 3674
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11716 2650 11744 3130
rect 12084 3126 12112 3334
rect 12912 3210 12940 3470
rect 13004 3398 13032 3878
rect 13084 3664 13136 3670
rect 13188 3618 13216 3878
rect 13136 3612 13216 3618
rect 13084 3606 13216 3612
rect 13096 3590 13216 3606
rect 13188 3398 13216 3590
rect 13556 3466 13584 4150
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13214 3292 13522 3301
rect 13214 3290 13220 3292
rect 13276 3290 13300 3292
rect 13356 3290 13380 3292
rect 13436 3290 13460 3292
rect 13516 3290 13522 3292
rect 13276 3238 13278 3290
rect 13458 3238 13460 3290
rect 13214 3236 13220 3238
rect 13276 3236 13300 3238
rect 13356 3236 13380 3238
rect 13436 3236 13460 3238
rect 13516 3236 13522 3238
rect 13214 3227 13522 3236
rect 12912 3182 13032 3210
rect 12072 3120 12124 3126
rect 12072 3062 12124 3068
rect 13004 2990 13032 3182
rect 13556 3058 13584 3402
rect 13648 3058 13676 4218
rect 13832 4162 13860 5170
rect 14016 5030 14044 5170
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 13924 4214 13952 4422
rect 14292 4214 14320 4422
rect 13740 4134 13860 4162
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 13740 3534 13768 4134
rect 13924 3942 13952 4150
rect 14476 4146 14504 4966
rect 14568 4826 14596 5102
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14660 4554 14688 5238
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 14752 4486 14780 5510
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14752 4146 14780 4422
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13924 3534 13952 3878
rect 14016 3738 14044 4014
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14292 3126 14320 3402
rect 14752 3194 14780 4082
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 4632 1170 4660 2314
rect 7214 2204 7522 2213
rect 7214 2202 7220 2204
rect 7276 2202 7300 2204
rect 7356 2202 7380 2204
rect 7436 2202 7460 2204
rect 7516 2202 7522 2204
rect 7276 2150 7278 2202
rect 7458 2150 7460 2202
rect 7214 2148 7220 2150
rect 7276 2148 7300 2150
rect 7356 2148 7380 2150
rect 7436 2148 7460 2150
rect 7516 2148 7522 2150
rect 7214 2139 7522 2148
rect 9784 1306 9812 2382
rect 13214 2204 13522 2213
rect 13214 2202 13220 2204
rect 13276 2202 13300 2204
rect 13356 2202 13380 2204
rect 13436 2202 13460 2204
rect 13516 2202 13522 2204
rect 13276 2150 13278 2202
rect 13458 2150 13460 2202
rect 13214 2148 13220 2150
rect 13276 2148 13300 2150
rect 13356 2148 13380 2150
rect 13436 2148 13460 2150
rect 13516 2148 13522 2150
rect 13214 2139 13522 2148
rect 4540 1142 4660 1170
rect 9692 1278 9812 1306
rect 4540 800 4568 1142
rect 9692 800 9720 1278
rect 14844 800 14872 9574
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15028 9042 15056 9318
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 15396 8838 15424 9318
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15120 7818 15148 8434
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15120 7410 15148 7754
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 15212 5370 15240 5578
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4162 15240 4422
rect 15120 4134 15240 4162
rect 15120 3126 15148 4134
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15304 3126 15332 3334
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15396 2650 15424 8774
rect 15488 8634 15516 9522
rect 15764 8974 15792 9930
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15856 9722 15884 9862
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 16132 9178 16160 10066
rect 16214 9276 16522 9285
rect 16214 9274 16220 9276
rect 16276 9274 16300 9276
rect 16356 9274 16380 9276
rect 16436 9274 16460 9276
rect 16516 9274 16522 9276
rect 16276 9222 16278 9274
rect 16458 9222 16460 9274
rect 16214 9220 16220 9222
rect 16276 9220 16300 9222
rect 16356 9220 16380 9222
rect 16436 9220 16460 9222
rect 16516 9220 16522 9222
rect 16214 9211 16522 9220
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 16500 8378 16528 8434
rect 15488 7546 15516 8366
rect 16500 8350 16620 8378
rect 16214 8188 16522 8197
rect 16214 8186 16220 8188
rect 16276 8186 16300 8188
rect 16356 8186 16380 8188
rect 16436 8186 16460 8188
rect 16516 8186 16522 8188
rect 16276 8134 16278 8186
rect 16458 8134 16460 8186
rect 16214 8132 16220 8134
rect 16276 8132 16300 8134
rect 16356 8132 16380 8134
rect 16436 8132 16460 8134
rect 16516 8132 16522 8134
rect 16214 8123 16522 8132
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15856 7546 15884 7686
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 16592 7410 16620 8350
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16214 7100 16522 7109
rect 16214 7098 16220 7100
rect 16276 7098 16300 7100
rect 16356 7098 16380 7100
rect 16436 7098 16460 7100
rect 16516 7098 16522 7100
rect 16276 7046 16278 7098
rect 16458 7046 16460 7098
rect 16214 7044 16220 7046
rect 16276 7044 16300 7046
rect 16356 7044 16380 7046
rect 16436 7044 16460 7046
rect 16516 7044 16522 7046
rect 16214 7035 16522 7044
rect 16592 7002 16620 7210
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 17130 6896 17186 6905
rect 17130 6831 17132 6840
rect 17184 6831 17186 6840
rect 17132 6802 17184 6808
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15672 5642 15700 6394
rect 16214 6012 16522 6021
rect 16214 6010 16220 6012
rect 16276 6010 16300 6012
rect 16356 6010 16380 6012
rect 16436 6010 16460 6012
rect 16516 6010 16522 6012
rect 16276 5958 16278 6010
rect 16458 5958 16460 6010
rect 16214 5956 16220 5958
rect 16276 5956 16300 5958
rect 16356 5956 16380 5958
rect 16436 5956 16460 5958
rect 16516 5956 16522 5958
rect 16214 5947 16522 5956
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 15672 5250 15700 5578
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 5302 16712 5510
rect 15580 5222 15700 5250
rect 16672 5296 16724 5302
rect 16672 5238 16724 5244
rect 15580 4486 15608 5222
rect 16214 4924 16522 4933
rect 16214 4922 16220 4924
rect 16276 4922 16300 4924
rect 16356 4922 16380 4924
rect 16436 4922 16460 4924
rect 16516 4922 16522 4924
rect 16276 4870 16278 4922
rect 16458 4870 16460 4922
rect 16214 4868 16220 4870
rect 16276 4868 16300 4870
rect 16356 4868 16380 4870
rect 16436 4868 16460 4870
rect 16516 4868 16522 4870
rect 16214 4859 16522 4868
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4214 15608 4422
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 16214 3836 16522 3845
rect 16214 3834 16220 3836
rect 16276 3834 16300 3836
rect 16356 3834 16380 3836
rect 16436 3834 16460 3836
rect 16516 3834 16522 3836
rect 16276 3782 16278 3834
rect 16458 3782 16460 3834
rect 16214 3780 16220 3782
rect 16276 3780 16300 3782
rect 16356 3780 16380 3782
rect 16436 3780 16460 3782
rect 16516 3780 16522 3782
rect 16214 3771 16522 3780
rect 16214 2748 16522 2757
rect 16214 2746 16220 2748
rect 16276 2746 16300 2748
rect 16356 2746 16380 2748
rect 16436 2746 16460 2748
rect 16516 2746 16522 2748
rect 16276 2694 16278 2746
rect 16458 2694 16460 2746
rect 16214 2692 16220 2694
rect 16276 2692 16300 2694
rect 16356 2692 16380 2694
rect 16436 2692 16460 2694
rect 16516 2692 16522 2694
rect 16214 2683 16522 2692
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17052 1465 17080 2382
rect 17038 1456 17094 1465
rect 17038 1391 17094 1400
rect 18 0 74 800
rect 4526 0 4582 800
rect 9678 0 9734 800
rect 14830 0 14886 800
<< via2 >>
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 10220 17978 10276 17980
rect 10300 17978 10356 17980
rect 10380 17978 10436 17980
rect 10460 17978 10516 17980
rect 10220 17926 10266 17978
rect 10266 17926 10276 17978
rect 10300 17926 10330 17978
rect 10330 17926 10342 17978
rect 10342 17926 10356 17978
rect 10380 17926 10394 17978
rect 10394 17926 10406 17978
rect 10406 17926 10436 17978
rect 10460 17926 10470 17978
rect 10470 17926 10516 17978
rect 10220 17924 10276 17926
rect 10300 17924 10356 17926
rect 10380 17924 10436 17926
rect 10460 17924 10516 17926
rect 7220 17434 7276 17436
rect 7300 17434 7356 17436
rect 7380 17434 7436 17436
rect 7460 17434 7516 17436
rect 7220 17382 7266 17434
rect 7266 17382 7276 17434
rect 7300 17382 7330 17434
rect 7330 17382 7342 17434
rect 7342 17382 7356 17434
rect 7380 17382 7394 17434
rect 7394 17382 7406 17434
rect 7406 17382 7436 17434
rect 7460 17382 7470 17434
rect 7470 17382 7516 17434
rect 7220 17380 7276 17382
rect 7300 17380 7356 17382
rect 7380 17380 7436 17382
rect 7460 17380 7516 17382
rect 16220 17978 16276 17980
rect 16300 17978 16356 17980
rect 16380 17978 16436 17980
rect 16460 17978 16516 17980
rect 16220 17926 16266 17978
rect 16266 17926 16276 17978
rect 16300 17926 16330 17978
rect 16330 17926 16342 17978
rect 16342 17926 16356 17978
rect 16380 17926 16394 17978
rect 16394 17926 16406 17978
rect 16406 17926 16436 17978
rect 16460 17926 16470 17978
rect 16470 17926 16516 17978
rect 16220 17924 16276 17926
rect 16300 17924 16356 17926
rect 16380 17924 16436 17926
rect 16460 17924 16516 17926
rect 17038 17740 17094 17776
rect 17038 17720 17040 17740
rect 17040 17720 17092 17740
rect 17092 17720 17094 17740
rect 13220 17434 13276 17436
rect 13300 17434 13356 17436
rect 13380 17434 13436 17436
rect 13460 17434 13516 17436
rect 13220 17382 13266 17434
rect 13266 17382 13276 17434
rect 13300 17382 13330 17434
rect 13330 17382 13342 17434
rect 13342 17382 13356 17434
rect 13380 17382 13394 17434
rect 13394 17382 13406 17434
rect 13406 17382 13436 17434
rect 13460 17382 13470 17434
rect 13470 17382 13516 17434
rect 13220 17380 13276 17382
rect 13300 17380 13356 17382
rect 13380 17380 13436 17382
rect 13460 17380 13516 17382
rect 10220 16890 10276 16892
rect 10300 16890 10356 16892
rect 10380 16890 10436 16892
rect 10460 16890 10516 16892
rect 10220 16838 10266 16890
rect 10266 16838 10276 16890
rect 10300 16838 10330 16890
rect 10330 16838 10342 16890
rect 10342 16838 10356 16890
rect 10380 16838 10394 16890
rect 10394 16838 10406 16890
rect 10406 16838 10436 16890
rect 10460 16838 10470 16890
rect 10470 16838 10516 16890
rect 10220 16836 10276 16838
rect 10300 16836 10356 16838
rect 10380 16836 10436 16838
rect 10460 16836 10516 16838
rect 938 15680 994 15736
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 938 10240 994 10296
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 7220 16346 7276 16348
rect 7300 16346 7356 16348
rect 7380 16346 7436 16348
rect 7460 16346 7516 16348
rect 7220 16294 7266 16346
rect 7266 16294 7276 16346
rect 7300 16294 7330 16346
rect 7330 16294 7342 16346
rect 7342 16294 7356 16346
rect 7380 16294 7394 16346
rect 7394 16294 7406 16346
rect 7406 16294 7436 16346
rect 7460 16294 7470 16346
rect 7470 16294 7516 16346
rect 7220 16292 7276 16294
rect 7300 16292 7356 16294
rect 7380 16292 7436 16294
rect 7460 16292 7516 16294
rect 10220 15802 10276 15804
rect 10300 15802 10356 15804
rect 10380 15802 10436 15804
rect 10460 15802 10516 15804
rect 10220 15750 10266 15802
rect 10266 15750 10276 15802
rect 10300 15750 10330 15802
rect 10330 15750 10342 15802
rect 10342 15750 10356 15802
rect 10380 15750 10394 15802
rect 10394 15750 10406 15802
rect 10406 15750 10436 15802
rect 10460 15750 10470 15802
rect 10470 15750 10516 15802
rect 10220 15748 10276 15750
rect 10300 15748 10356 15750
rect 10380 15748 10436 15750
rect 10460 15748 10516 15750
rect 16220 16890 16276 16892
rect 16300 16890 16356 16892
rect 16380 16890 16436 16892
rect 16460 16890 16516 16892
rect 16220 16838 16266 16890
rect 16266 16838 16276 16890
rect 16300 16838 16330 16890
rect 16330 16838 16342 16890
rect 16342 16838 16356 16890
rect 16380 16838 16394 16890
rect 16394 16838 16406 16890
rect 16406 16838 16436 16890
rect 16460 16838 16470 16890
rect 16470 16838 16516 16890
rect 16220 16836 16276 16838
rect 16300 16836 16356 16838
rect 16380 16836 16436 16838
rect 16460 16836 16516 16838
rect 13220 16346 13276 16348
rect 13300 16346 13356 16348
rect 13380 16346 13436 16348
rect 13460 16346 13516 16348
rect 13220 16294 13266 16346
rect 13266 16294 13276 16346
rect 13300 16294 13330 16346
rect 13330 16294 13342 16346
rect 13342 16294 13356 16346
rect 13380 16294 13394 16346
rect 13394 16294 13406 16346
rect 13406 16294 13436 16346
rect 13460 16294 13470 16346
rect 13470 16294 13516 16346
rect 13220 16292 13276 16294
rect 13300 16292 13356 16294
rect 13380 16292 13436 16294
rect 13460 16292 13516 16294
rect 7220 15258 7276 15260
rect 7300 15258 7356 15260
rect 7380 15258 7436 15260
rect 7460 15258 7516 15260
rect 7220 15206 7266 15258
rect 7266 15206 7276 15258
rect 7300 15206 7330 15258
rect 7330 15206 7342 15258
rect 7342 15206 7356 15258
rect 7380 15206 7394 15258
rect 7394 15206 7406 15258
rect 7406 15206 7436 15258
rect 7460 15206 7470 15258
rect 7470 15206 7516 15258
rect 7220 15204 7276 15206
rect 7300 15204 7356 15206
rect 7380 15204 7436 15206
rect 7460 15204 7516 15206
rect 7220 14170 7276 14172
rect 7300 14170 7356 14172
rect 7380 14170 7436 14172
rect 7460 14170 7516 14172
rect 7220 14118 7266 14170
rect 7266 14118 7276 14170
rect 7300 14118 7330 14170
rect 7330 14118 7342 14170
rect 7342 14118 7356 14170
rect 7380 14118 7394 14170
rect 7394 14118 7406 14170
rect 7406 14118 7436 14170
rect 7460 14118 7470 14170
rect 7470 14118 7516 14170
rect 7220 14116 7276 14118
rect 7300 14116 7356 14118
rect 7380 14116 7436 14118
rect 7460 14116 7516 14118
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 7220 13082 7276 13084
rect 7300 13082 7356 13084
rect 7380 13082 7436 13084
rect 7460 13082 7516 13084
rect 7220 13030 7266 13082
rect 7266 13030 7276 13082
rect 7300 13030 7330 13082
rect 7330 13030 7342 13082
rect 7342 13030 7356 13082
rect 7380 13030 7394 13082
rect 7394 13030 7406 13082
rect 7406 13030 7436 13082
rect 7460 13030 7470 13082
rect 7470 13030 7516 13082
rect 7220 13028 7276 13030
rect 7300 13028 7356 13030
rect 7380 13028 7436 13030
rect 7460 13028 7516 13030
rect 7220 11994 7276 11996
rect 7300 11994 7356 11996
rect 7380 11994 7436 11996
rect 7460 11994 7516 11996
rect 7220 11942 7266 11994
rect 7266 11942 7276 11994
rect 7300 11942 7330 11994
rect 7330 11942 7342 11994
rect 7342 11942 7356 11994
rect 7380 11942 7394 11994
rect 7394 11942 7406 11994
rect 7406 11942 7436 11994
rect 7460 11942 7470 11994
rect 7470 11942 7516 11994
rect 7220 11940 7276 11942
rect 7300 11940 7356 11942
rect 7380 11940 7436 11942
rect 7460 11940 7516 11942
rect 7220 10906 7276 10908
rect 7300 10906 7356 10908
rect 7380 10906 7436 10908
rect 7460 10906 7516 10908
rect 7220 10854 7266 10906
rect 7266 10854 7276 10906
rect 7300 10854 7330 10906
rect 7330 10854 7342 10906
rect 7342 10854 7356 10906
rect 7380 10854 7394 10906
rect 7394 10854 7406 10906
rect 7406 10854 7436 10906
rect 7460 10854 7470 10906
rect 7470 10854 7516 10906
rect 7220 10852 7276 10854
rect 7300 10852 7356 10854
rect 7380 10852 7436 10854
rect 7460 10852 7516 10854
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 7220 9818 7276 9820
rect 7300 9818 7356 9820
rect 7380 9818 7436 9820
rect 7460 9818 7516 9820
rect 7220 9766 7266 9818
rect 7266 9766 7276 9818
rect 7300 9766 7330 9818
rect 7330 9766 7342 9818
rect 7342 9766 7356 9818
rect 7380 9766 7394 9818
rect 7394 9766 7406 9818
rect 7406 9766 7436 9818
rect 7460 9766 7470 9818
rect 7470 9766 7516 9818
rect 7220 9764 7276 9766
rect 7300 9764 7356 9766
rect 7380 9764 7436 9766
rect 7460 9764 7516 9766
rect 7220 8730 7276 8732
rect 7300 8730 7356 8732
rect 7380 8730 7436 8732
rect 7460 8730 7516 8732
rect 7220 8678 7266 8730
rect 7266 8678 7276 8730
rect 7300 8678 7330 8730
rect 7330 8678 7342 8730
rect 7342 8678 7356 8730
rect 7380 8678 7394 8730
rect 7394 8678 7406 8730
rect 7406 8678 7436 8730
rect 7460 8678 7470 8730
rect 7470 8678 7516 8730
rect 7220 8676 7276 8678
rect 7300 8676 7356 8678
rect 7380 8676 7436 8678
rect 7460 8676 7516 8678
rect 10220 14714 10276 14716
rect 10300 14714 10356 14716
rect 10380 14714 10436 14716
rect 10460 14714 10516 14716
rect 10220 14662 10266 14714
rect 10266 14662 10276 14714
rect 10300 14662 10330 14714
rect 10330 14662 10342 14714
rect 10342 14662 10356 14714
rect 10380 14662 10394 14714
rect 10394 14662 10406 14714
rect 10406 14662 10436 14714
rect 10460 14662 10470 14714
rect 10470 14662 10516 14714
rect 10220 14660 10276 14662
rect 10300 14660 10356 14662
rect 10380 14660 10436 14662
rect 10460 14660 10516 14662
rect 10220 13626 10276 13628
rect 10300 13626 10356 13628
rect 10380 13626 10436 13628
rect 10460 13626 10516 13628
rect 10220 13574 10266 13626
rect 10266 13574 10276 13626
rect 10300 13574 10330 13626
rect 10330 13574 10342 13626
rect 10342 13574 10356 13626
rect 10380 13574 10394 13626
rect 10394 13574 10406 13626
rect 10406 13574 10436 13626
rect 10460 13574 10470 13626
rect 10470 13574 10516 13626
rect 10220 13572 10276 13574
rect 10300 13572 10356 13574
rect 10380 13572 10436 13574
rect 10460 13572 10516 13574
rect 10220 12538 10276 12540
rect 10300 12538 10356 12540
rect 10380 12538 10436 12540
rect 10460 12538 10516 12540
rect 10220 12486 10266 12538
rect 10266 12486 10276 12538
rect 10300 12486 10330 12538
rect 10330 12486 10342 12538
rect 10342 12486 10356 12538
rect 10380 12486 10394 12538
rect 10394 12486 10406 12538
rect 10406 12486 10436 12538
rect 10460 12486 10470 12538
rect 10470 12486 10516 12538
rect 10220 12484 10276 12486
rect 10300 12484 10356 12486
rect 10380 12484 10436 12486
rect 10460 12484 10516 12486
rect 10220 11450 10276 11452
rect 10300 11450 10356 11452
rect 10380 11450 10436 11452
rect 10460 11450 10516 11452
rect 10220 11398 10266 11450
rect 10266 11398 10276 11450
rect 10300 11398 10330 11450
rect 10330 11398 10342 11450
rect 10342 11398 10356 11450
rect 10380 11398 10394 11450
rect 10394 11398 10406 11450
rect 10406 11398 10436 11450
rect 10460 11398 10470 11450
rect 10470 11398 10516 11450
rect 10220 11396 10276 11398
rect 10300 11396 10356 11398
rect 10380 11396 10436 11398
rect 10460 11396 10516 11398
rect 10220 10362 10276 10364
rect 10300 10362 10356 10364
rect 10380 10362 10436 10364
rect 10460 10362 10516 10364
rect 10220 10310 10266 10362
rect 10266 10310 10276 10362
rect 10300 10310 10330 10362
rect 10330 10310 10342 10362
rect 10342 10310 10356 10362
rect 10380 10310 10394 10362
rect 10394 10310 10406 10362
rect 10406 10310 10436 10362
rect 10460 10310 10470 10362
rect 10470 10310 10516 10362
rect 10220 10308 10276 10310
rect 10300 10308 10356 10310
rect 10380 10308 10436 10310
rect 10460 10308 10516 10310
rect 10220 9274 10276 9276
rect 10300 9274 10356 9276
rect 10380 9274 10436 9276
rect 10460 9274 10516 9276
rect 10220 9222 10266 9274
rect 10266 9222 10276 9274
rect 10300 9222 10330 9274
rect 10330 9222 10342 9274
rect 10342 9222 10356 9274
rect 10380 9222 10394 9274
rect 10394 9222 10406 9274
rect 10406 9222 10436 9274
rect 10460 9222 10470 9274
rect 10470 9222 10516 9274
rect 10220 9220 10276 9222
rect 10300 9220 10356 9222
rect 10380 9220 10436 9222
rect 10460 9220 10516 9222
rect 10220 8186 10276 8188
rect 10300 8186 10356 8188
rect 10380 8186 10436 8188
rect 10460 8186 10516 8188
rect 10220 8134 10266 8186
rect 10266 8134 10276 8186
rect 10300 8134 10330 8186
rect 10330 8134 10342 8186
rect 10342 8134 10356 8186
rect 10380 8134 10394 8186
rect 10394 8134 10406 8186
rect 10406 8134 10436 8186
rect 10460 8134 10470 8186
rect 10470 8134 10516 8186
rect 10220 8132 10276 8134
rect 10300 8132 10356 8134
rect 10380 8132 10436 8134
rect 10460 8132 10516 8134
rect 7220 7642 7276 7644
rect 7300 7642 7356 7644
rect 7380 7642 7436 7644
rect 7460 7642 7516 7644
rect 7220 7590 7266 7642
rect 7266 7590 7276 7642
rect 7300 7590 7330 7642
rect 7330 7590 7342 7642
rect 7342 7590 7356 7642
rect 7380 7590 7394 7642
rect 7394 7590 7406 7642
rect 7406 7590 7436 7642
rect 7460 7590 7470 7642
rect 7470 7590 7516 7642
rect 7220 7588 7276 7590
rect 7300 7588 7356 7590
rect 7380 7588 7436 7590
rect 7460 7588 7516 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 938 4800 994 4856
rect 7220 6554 7276 6556
rect 7300 6554 7356 6556
rect 7380 6554 7436 6556
rect 7460 6554 7516 6556
rect 7220 6502 7266 6554
rect 7266 6502 7276 6554
rect 7300 6502 7330 6554
rect 7330 6502 7342 6554
rect 7342 6502 7356 6554
rect 7380 6502 7394 6554
rect 7394 6502 7406 6554
rect 7406 6502 7436 6554
rect 7460 6502 7470 6554
rect 7470 6502 7516 6554
rect 7220 6500 7276 6502
rect 7300 6500 7356 6502
rect 7380 6500 7436 6502
rect 7460 6500 7516 6502
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 7220 5466 7276 5468
rect 7300 5466 7356 5468
rect 7380 5466 7436 5468
rect 7460 5466 7516 5468
rect 7220 5414 7266 5466
rect 7266 5414 7276 5466
rect 7300 5414 7330 5466
rect 7330 5414 7342 5466
rect 7342 5414 7356 5466
rect 7380 5414 7394 5466
rect 7394 5414 7406 5466
rect 7406 5414 7436 5466
rect 7460 5414 7470 5466
rect 7470 5414 7516 5466
rect 7220 5412 7276 5414
rect 7300 5412 7356 5414
rect 7380 5412 7436 5414
rect 7460 5412 7516 5414
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 7220 4378 7276 4380
rect 7300 4378 7356 4380
rect 7380 4378 7436 4380
rect 7460 4378 7516 4380
rect 7220 4326 7266 4378
rect 7266 4326 7276 4378
rect 7300 4326 7330 4378
rect 7330 4326 7342 4378
rect 7342 4326 7356 4378
rect 7380 4326 7394 4378
rect 7394 4326 7406 4378
rect 7406 4326 7436 4378
rect 7460 4326 7470 4378
rect 7470 4326 7516 4378
rect 7220 4324 7276 4326
rect 7300 4324 7356 4326
rect 7380 4324 7436 4326
rect 7460 4324 7516 4326
rect 10220 7098 10276 7100
rect 10300 7098 10356 7100
rect 10380 7098 10436 7100
rect 10460 7098 10516 7100
rect 10220 7046 10266 7098
rect 10266 7046 10276 7098
rect 10300 7046 10330 7098
rect 10330 7046 10342 7098
rect 10342 7046 10356 7098
rect 10380 7046 10394 7098
rect 10394 7046 10406 7098
rect 10406 7046 10436 7098
rect 10460 7046 10470 7098
rect 10470 7046 10516 7098
rect 10220 7044 10276 7046
rect 10300 7044 10356 7046
rect 10380 7044 10436 7046
rect 10460 7044 10516 7046
rect 10220 6010 10276 6012
rect 10300 6010 10356 6012
rect 10380 6010 10436 6012
rect 10460 6010 10516 6012
rect 10220 5958 10266 6010
rect 10266 5958 10276 6010
rect 10300 5958 10330 6010
rect 10330 5958 10342 6010
rect 10342 5958 10356 6010
rect 10380 5958 10394 6010
rect 10394 5958 10406 6010
rect 10406 5958 10436 6010
rect 10460 5958 10470 6010
rect 10470 5958 10516 6010
rect 10220 5956 10276 5958
rect 10300 5956 10356 5958
rect 10380 5956 10436 5958
rect 10460 5956 10516 5958
rect 10220 4922 10276 4924
rect 10300 4922 10356 4924
rect 10380 4922 10436 4924
rect 10460 4922 10516 4924
rect 10220 4870 10266 4922
rect 10266 4870 10276 4922
rect 10300 4870 10330 4922
rect 10330 4870 10342 4922
rect 10342 4870 10356 4922
rect 10380 4870 10394 4922
rect 10394 4870 10406 4922
rect 10406 4870 10436 4922
rect 10460 4870 10470 4922
rect 10470 4870 10516 4922
rect 10220 4868 10276 4870
rect 10300 4868 10356 4870
rect 10380 4868 10436 4870
rect 10460 4868 10516 4870
rect 7220 3290 7276 3292
rect 7300 3290 7356 3292
rect 7380 3290 7436 3292
rect 7460 3290 7516 3292
rect 7220 3238 7266 3290
rect 7266 3238 7276 3290
rect 7300 3238 7330 3290
rect 7330 3238 7342 3290
rect 7342 3238 7356 3290
rect 7380 3238 7394 3290
rect 7394 3238 7406 3290
rect 7406 3238 7436 3290
rect 7460 3238 7470 3290
rect 7470 3238 7516 3290
rect 7220 3236 7276 3238
rect 7300 3236 7356 3238
rect 7380 3236 7436 3238
rect 7460 3236 7516 3238
rect 10220 3834 10276 3836
rect 10300 3834 10356 3836
rect 10380 3834 10436 3836
rect 10460 3834 10516 3836
rect 10220 3782 10266 3834
rect 10266 3782 10276 3834
rect 10300 3782 10330 3834
rect 10330 3782 10342 3834
rect 10342 3782 10356 3834
rect 10380 3782 10394 3834
rect 10394 3782 10406 3834
rect 10406 3782 10436 3834
rect 10460 3782 10470 3834
rect 10470 3782 10516 3834
rect 10220 3780 10276 3782
rect 10300 3780 10356 3782
rect 10380 3780 10436 3782
rect 10460 3780 10516 3782
rect 10220 2746 10276 2748
rect 10300 2746 10356 2748
rect 10380 2746 10436 2748
rect 10460 2746 10516 2748
rect 10220 2694 10266 2746
rect 10266 2694 10276 2746
rect 10300 2694 10330 2746
rect 10330 2694 10342 2746
rect 10342 2694 10356 2746
rect 10380 2694 10394 2746
rect 10394 2694 10406 2746
rect 10406 2694 10436 2746
rect 10460 2694 10470 2746
rect 10470 2694 10516 2746
rect 10220 2692 10276 2694
rect 10300 2692 10356 2694
rect 10380 2692 10436 2694
rect 10460 2692 10516 2694
rect 13220 15258 13276 15260
rect 13300 15258 13356 15260
rect 13380 15258 13436 15260
rect 13460 15258 13516 15260
rect 13220 15206 13266 15258
rect 13266 15206 13276 15258
rect 13300 15206 13330 15258
rect 13330 15206 13342 15258
rect 13342 15206 13356 15258
rect 13380 15206 13394 15258
rect 13394 15206 13406 15258
rect 13406 15206 13436 15258
rect 13460 15206 13470 15258
rect 13470 15206 13516 15258
rect 13220 15204 13276 15206
rect 13300 15204 13356 15206
rect 13380 15204 13436 15206
rect 13460 15204 13516 15206
rect 16220 15802 16276 15804
rect 16300 15802 16356 15804
rect 16380 15802 16436 15804
rect 16460 15802 16516 15804
rect 16220 15750 16266 15802
rect 16266 15750 16276 15802
rect 16300 15750 16330 15802
rect 16330 15750 16342 15802
rect 16342 15750 16356 15802
rect 16380 15750 16394 15802
rect 16394 15750 16406 15802
rect 16406 15750 16436 15802
rect 16460 15750 16470 15802
rect 16470 15750 16516 15802
rect 16220 15748 16276 15750
rect 16300 15748 16356 15750
rect 16380 15748 16436 15750
rect 16460 15748 16516 15750
rect 13220 14170 13276 14172
rect 13300 14170 13356 14172
rect 13380 14170 13436 14172
rect 13460 14170 13516 14172
rect 13220 14118 13266 14170
rect 13266 14118 13276 14170
rect 13300 14118 13330 14170
rect 13330 14118 13342 14170
rect 13342 14118 13356 14170
rect 13380 14118 13394 14170
rect 13394 14118 13406 14170
rect 13406 14118 13436 14170
rect 13460 14118 13470 14170
rect 13470 14118 13516 14170
rect 13220 14116 13276 14118
rect 13300 14116 13356 14118
rect 13380 14116 13436 14118
rect 13460 14116 13516 14118
rect 13220 13082 13276 13084
rect 13300 13082 13356 13084
rect 13380 13082 13436 13084
rect 13460 13082 13516 13084
rect 13220 13030 13266 13082
rect 13266 13030 13276 13082
rect 13300 13030 13330 13082
rect 13330 13030 13342 13082
rect 13342 13030 13356 13082
rect 13380 13030 13394 13082
rect 13394 13030 13406 13082
rect 13406 13030 13436 13082
rect 13460 13030 13470 13082
rect 13470 13030 13516 13082
rect 13220 13028 13276 13030
rect 13300 13028 13356 13030
rect 13380 13028 13436 13030
rect 13460 13028 13516 13030
rect 13220 11994 13276 11996
rect 13300 11994 13356 11996
rect 13380 11994 13436 11996
rect 13460 11994 13516 11996
rect 13220 11942 13266 11994
rect 13266 11942 13276 11994
rect 13300 11942 13330 11994
rect 13330 11942 13342 11994
rect 13342 11942 13356 11994
rect 13380 11942 13394 11994
rect 13394 11942 13406 11994
rect 13406 11942 13436 11994
rect 13460 11942 13470 11994
rect 13470 11942 13516 11994
rect 13220 11940 13276 11942
rect 13300 11940 13356 11942
rect 13380 11940 13436 11942
rect 13460 11940 13516 11942
rect 13220 10906 13276 10908
rect 13300 10906 13356 10908
rect 13380 10906 13436 10908
rect 13460 10906 13516 10908
rect 13220 10854 13266 10906
rect 13266 10854 13276 10906
rect 13300 10854 13330 10906
rect 13330 10854 13342 10906
rect 13342 10854 13356 10906
rect 13380 10854 13394 10906
rect 13394 10854 13406 10906
rect 13406 10854 13436 10906
rect 13460 10854 13470 10906
rect 13470 10854 13516 10906
rect 13220 10852 13276 10854
rect 13300 10852 13356 10854
rect 13380 10852 13436 10854
rect 13460 10852 13516 10854
rect 13220 9818 13276 9820
rect 13300 9818 13356 9820
rect 13380 9818 13436 9820
rect 13460 9818 13516 9820
rect 13220 9766 13266 9818
rect 13266 9766 13276 9818
rect 13300 9766 13330 9818
rect 13330 9766 13342 9818
rect 13342 9766 13356 9818
rect 13380 9766 13394 9818
rect 13394 9766 13406 9818
rect 13406 9766 13436 9818
rect 13460 9766 13470 9818
rect 13470 9766 13516 9818
rect 13220 9764 13276 9766
rect 13300 9764 13356 9766
rect 13380 9764 13436 9766
rect 13460 9764 13516 9766
rect 16220 14714 16276 14716
rect 16300 14714 16356 14716
rect 16380 14714 16436 14716
rect 16460 14714 16516 14716
rect 16220 14662 16266 14714
rect 16266 14662 16276 14714
rect 16300 14662 16330 14714
rect 16330 14662 16342 14714
rect 16342 14662 16356 14714
rect 16380 14662 16394 14714
rect 16394 14662 16406 14714
rect 16406 14662 16436 14714
rect 16460 14662 16470 14714
rect 16470 14662 16516 14714
rect 16220 14660 16276 14662
rect 16300 14660 16356 14662
rect 16380 14660 16436 14662
rect 16460 14660 16516 14662
rect 16220 13626 16276 13628
rect 16300 13626 16356 13628
rect 16380 13626 16436 13628
rect 16460 13626 16516 13628
rect 16220 13574 16266 13626
rect 16266 13574 16276 13626
rect 16300 13574 16330 13626
rect 16330 13574 16342 13626
rect 16342 13574 16356 13626
rect 16380 13574 16394 13626
rect 16394 13574 16406 13626
rect 16406 13574 16436 13626
rect 16460 13574 16470 13626
rect 16470 13574 16516 13626
rect 16220 13572 16276 13574
rect 16300 13572 16356 13574
rect 16380 13572 16436 13574
rect 16460 13572 16516 13574
rect 16220 12538 16276 12540
rect 16300 12538 16356 12540
rect 16380 12538 16436 12540
rect 16460 12538 16516 12540
rect 16220 12486 16266 12538
rect 16266 12486 16276 12538
rect 16300 12486 16330 12538
rect 16330 12486 16342 12538
rect 16342 12486 16356 12538
rect 16380 12486 16394 12538
rect 16394 12486 16406 12538
rect 16406 12486 16436 12538
rect 16460 12486 16470 12538
rect 16470 12486 16516 12538
rect 16220 12484 16276 12486
rect 16300 12484 16356 12486
rect 16380 12484 16436 12486
rect 16460 12484 16516 12486
rect 16118 12280 16174 12336
rect 16220 11450 16276 11452
rect 16300 11450 16356 11452
rect 16380 11450 16436 11452
rect 16460 11450 16516 11452
rect 16220 11398 16266 11450
rect 16266 11398 16276 11450
rect 16300 11398 16330 11450
rect 16330 11398 16342 11450
rect 16342 11398 16356 11450
rect 16380 11398 16394 11450
rect 16394 11398 16406 11450
rect 16406 11398 16436 11450
rect 16460 11398 16470 11450
rect 16470 11398 16516 11450
rect 16220 11396 16276 11398
rect 16300 11396 16356 11398
rect 16380 11396 16436 11398
rect 16460 11396 16516 11398
rect 16220 10362 16276 10364
rect 16300 10362 16356 10364
rect 16380 10362 16436 10364
rect 16460 10362 16516 10364
rect 16220 10310 16266 10362
rect 16266 10310 16276 10362
rect 16300 10310 16330 10362
rect 16330 10310 16342 10362
rect 16342 10310 16356 10362
rect 16380 10310 16394 10362
rect 16394 10310 16406 10362
rect 16406 10310 16436 10362
rect 16460 10310 16470 10362
rect 16470 10310 16516 10362
rect 16220 10308 16276 10310
rect 16300 10308 16356 10310
rect 16380 10308 16436 10310
rect 16460 10308 16516 10310
rect 13220 8730 13276 8732
rect 13300 8730 13356 8732
rect 13380 8730 13436 8732
rect 13460 8730 13516 8732
rect 13220 8678 13266 8730
rect 13266 8678 13276 8730
rect 13300 8678 13330 8730
rect 13330 8678 13342 8730
rect 13342 8678 13356 8730
rect 13380 8678 13394 8730
rect 13394 8678 13406 8730
rect 13406 8678 13436 8730
rect 13460 8678 13470 8730
rect 13470 8678 13516 8730
rect 13220 8676 13276 8678
rect 13300 8676 13356 8678
rect 13380 8676 13436 8678
rect 13460 8676 13516 8678
rect 13220 7642 13276 7644
rect 13300 7642 13356 7644
rect 13380 7642 13436 7644
rect 13460 7642 13516 7644
rect 13220 7590 13266 7642
rect 13266 7590 13276 7642
rect 13300 7590 13330 7642
rect 13330 7590 13342 7642
rect 13342 7590 13356 7642
rect 13380 7590 13394 7642
rect 13394 7590 13406 7642
rect 13406 7590 13436 7642
rect 13460 7590 13470 7642
rect 13470 7590 13516 7642
rect 13220 7588 13276 7590
rect 13300 7588 13356 7590
rect 13380 7588 13436 7590
rect 13460 7588 13516 7590
rect 13220 6554 13276 6556
rect 13300 6554 13356 6556
rect 13380 6554 13436 6556
rect 13460 6554 13516 6556
rect 13220 6502 13266 6554
rect 13266 6502 13276 6554
rect 13300 6502 13330 6554
rect 13330 6502 13342 6554
rect 13342 6502 13356 6554
rect 13380 6502 13394 6554
rect 13394 6502 13406 6554
rect 13406 6502 13436 6554
rect 13460 6502 13470 6554
rect 13470 6502 13516 6554
rect 13220 6500 13276 6502
rect 13300 6500 13356 6502
rect 13380 6500 13436 6502
rect 13460 6500 13516 6502
rect 13220 5466 13276 5468
rect 13300 5466 13356 5468
rect 13380 5466 13436 5468
rect 13460 5466 13516 5468
rect 13220 5414 13266 5466
rect 13266 5414 13276 5466
rect 13300 5414 13330 5466
rect 13330 5414 13342 5466
rect 13342 5414 13356 5466
rect 13380 5414 13394 5466
rect 13394 5414 13406 5466
rect 13406 5414 13436 5466
rect 13460 5414 13470 5466
rect 13470 5414 13516 5466
rect 13220 5412 13276 5414
rect 13300 5412 13356 5414
rect 13380 5412 13436 5414
rect 13460 5412 13516 5414
rect 13220 4378 13276 4380
rect 13300 4378 13356 4380
rect 13380 4378 13436 4380
rect 13460 4378 13516 4380
rect 13220 4326 13266 4378
rect 13266 4326 13276 4378
rect 13300 4326 13330 4378
rect 13330 4326 13342 4378
rect 13342 4326 13356 4378
rect 13380 4326 13394 4378
rect 13394 4326 13406 4378
rect 13406 4326 13436 4378
rect 13460 4326 13470 4378
rect 13470 4326 13516 4378
rect 13220 4324 13276 4326
rect 13300 4324 13356 4326
rect 13380 4324 13436 4326
rect 13460 4324 13516 4326
rect 13220 3290 13276 3292
rect 13300 3290 13356 3292
rect 13380 3290 13436 3292
rect 13460 3290 13516 3292
rect 13220 3238 13266 3290
rect 13266 3238 13276 3290
rect 13300 3238 13330 3290
rect 13330 3238 13342 3290
rect 13342 3238 13356 3290
rect 13380 3238 13394 3290
rect 13394 3238 13406 3290
rect 13406 3238 13436 3290
rect 13460 3238 13470 3290
rect 13470 3238 13516 3290
rect 13220 3236 13276 3238
rect 13300 3236 13356 3238
rect 13380 3236 13436 3238
rect 13460 3236 13516 3238
rect 7220 2202 7276 2204
rect 7300 2202 7356 2204
rect 7380 2202 7436 2204
rect 7460 2202 7516 2204
rect 7220 2150 7266 2202
rect 7266 2150 7276 2202
rect 7300 2150 7330 2202
rect 7330 2150 7342 2202
rect 7342 2150 7356 2202
rect 7380 2150 7394 2202
rect 7394 2150 7406 2202
rect 7406 2150 7436 2202
rect 7460 2150 7470 2202
rect 7470 2150 7516 2202
rect 7220 2148 7276 2150
rect 7300 2148 7356 2150
rect 7380 2148 7436 2150
rect 7460 2148 7516 2150
rect 13220 2202 13276 2204
rect 13300 2202 13356 2204
rect 13380 2202 13436 2204
rect 13460 2202 13516 2204
rect 13220 2150 13266 2202
rect 13266 2150 13276 2202
rect 13300 2150 13330 2202
rect 13330 2150 13342 2202
rect 13342 2150 13356 2202
rect 13380 2150 13394 2202
rect 13394 2150 13406 2202
rect 13406 2150 13436 2202
rect 13460 2150 13470 2202
rect 13470 2150 13516 2202
rect 13220 2148 13276 2150
rect 13300 2148 13356 2150
rect 13380 2148 13436 2150
rect 13460 2148 13516 2150
rect 16220 9274 16276 9276
rect 16300 9274 16356 9276
rect 16380 9274 16436 9276
rect 16460 9274 16516 9276
rect 16220 9222 16266 9274
rect 16266 9222 16276 9274
rect 16300 9222 16330 9274
rect 16330 9222 16342 9274
rect 16342 9222 16356 9274
rect 16380 9222 16394 9274
rect 16394 9222 16406 9274
rect 16406 9222 16436 9274
rect 16460 9222 16470 9274
rect 16470 9222 16516 9274
rect 16220 9220 16276 9222
rect 16300 9220 16356 9222
rect 16380 9220 16436 9222
rect 16460 9220 16516 9222
rect 16220 8186 16276 8188
rect 16300 8186 16356 8188
rect 16380 8186 16436 8188
rect 16460 8186 16516 8188
rect 16220 8134 16266 8186
rect 16266 8134 16276 8186
rect 16300 8134 16330 8186
rect 16330 8134 16342 8186
rect 16342 8134 16356 8186
rect 16380 8134 16394 8186
rect 16394 8134 16406 8186
rect 16406 8134 16436 8186
rect 16460 8134 16470 8186
rect 16470 8134 16516 8186
rect 16220 8132 16276 8134
rect 16300 8132 16356 8134
rect 16380 8132 16436 8134
rect 16460 8132 16516 8134
rect 16220 7098 16276 7100
rect 16300 7098 16356 7100
rect 16380 7098 16436 7100
rect 16460 7098 16516 7100
rect 16220 7046 16266 7098
rect 16266 7046 16276 7098
rect 16300 7046 16330 7098
rect 16330 7046 16342 7098
rect 16342 7046 16356 7098
rect 16380 7046 16394 7098
rect 16394 7046 16406 7098
rect 16406 7046 16436 7098
rect 16460 7046 16470 7098
rect 16470 7046 16516 7098
rect 16220 7044 16276 7046
rect 16300 7044 16356 7046
rect 16380 7044 16436 7046
rect 16460 7044 16516 7046
rect 17130 6860 17186 6896
rect 17130 6840 17132 6860
rect 17132 6840 17184 6860
rect 17184 6840 17186 6860
rect 16220 6010 16276 6012
rect 16300 6010 16356 6012
rect 16380 6010 16436 6012
rect 16460 6010 16516 6012
rect 16220 5958 16266 6010
rect 16266 5958 16276 6010
rect 16300 5958 16330 6010
rect 16330 5958 16342 6010
rect 16342 5958 16356 6010
rect 16380 5958 16394 6010
rect 16394 5958 16406 6010
rect 16406 5958 16436 6010
rect 16460 5958 16470 6010
rect 16470 5958 16516 6010
rect 16220 5956 16276 5958
rect 16300 5956 16356 5958
rect 16380 5956 16436 5958
rect 16460 5956 16516 5958
rect 16220 4922 16276 4924
rect 16300 4922 16356 4924
rect 16380 4922 16436 4924
rect 16460 4922 16516 4924
rect 16220 4870 16266 4922
rect 16266 4870 16276 4922
rect 16300 4870 16330 4922
rect 16330 4870 16342 4922
rect 16342 4870 16356 4922
rect 16380 4870 16394 4922
rect 16394 4870 16406 4922
rect 16406 4870 16436 4922
rect 16460 4870 16470 4922
rect 16470 4870 16516 4922
rect 16220 4868 16276 4870
rect 16300 4868 16356 4870
rect 16380 4868 16436 4870
rect 16460 4868 16516 4870
rect 16220 3834 16276 3836
rect 16300 3834 16356 3836
rect 16380 3834 16436 3836
rect 16460 3834 16516 3836
rect 16220 3782 16266 3834
rect 16266 3782 16276 3834
rect 16300 3782 16330 3834
rect 16330 3782 16342 3834
rect 16342 3782 16356 3834
rect 16380 3782 16394 3834
rect 16394 3782 16406 3834
rect 16406 3782 16436 3834
rect 16460 3782 16470 3834
rect 16470 3782 16516 3834
rect 16220 3780 16276 3782
rect 16300 3780 16356 3782
rect 16380 3780 16436 3782
rect 16460 3780 16516 3782
rect 16220 2746 16276 2748
rect 16300 2746 16356 2748
rect 16380 2746 16436 2748
rect 16460 2746 16516 2748
rect 16220 2694 16266 2746
rect 16266 2694 16276 2746
rect 16300 2694 16330 2746
rect 16330 2694 16342 2746
rect 16342 2694 16356 2746
rect 16380 2694 16394 2746
rect 16394 2694 16406 2746
rect 16406 2694 16436 2746
rect 16460 2694 16470 2746
rect 16470 2694 16516 2746
rect 16220 2692 16276 2694
rect 16300 2692 16356 2694
rect 16380 2692 16436 2694
rect 16460 2692 16516 2694
rect 17038 1400 17094 1456
<< metal3 >>
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 10210 17984 10526 17985
rect 10210 17920 10216 17984
rect 10280 17920 10296 17984
rect 10360 17920 10376 17984
rect 10440 17920 10456 17984
rect 10520 17920 10526 17984
rect 10210 17919 10526 17920
rect 16210 17984 16526 17985
rect 16210 17920 16216 17984
rect 16280 17920 16296 17984
rect 16360 17920 16376 17984
rect 16440 17920 16456 17984
rect 16520 17920 16526 17984
rect 16210 17919 16526 17920
rect 17033 17778 17099 17781
rect 17506 17778 18306 17808
rect 17033 17776 18306 17778
rect 17033 17720 17038 17776
rect 17094 17720 18306 17776
rect 17033 17718 18306 17720
rect 17033 17715 17099 17718
rect 17506 17688 18306 17718
rect 7210 17440 7526 17441
rect 7210 17376 7216 17440
rect 7280 17376 7296 17440
rect 7360 17376 7376 17440
rect 7440 17376 7456 17440
rect 7520 17376 7526 17440
rect 7210 17375 7526 17376
rect 13210 17440 13526 17441
rect 13210 17376 13216 17440
rect 13280 17376 13296 17440
rect 13360 17376 13376 17440
rect 13440 17376 13456 17440
rect 13520 17376 13526 17440
rect 13210 17375 13526 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 10210 16896 10526 16897
rect 10210 16832 10216 16896
rect 10280 16832 10296 16896
rect 10360 16832 10376 16896
rect 10440 16832 10456 16896
rect 10520 16832 10526 16896
rect 10210 16831 10526 16832
rect 16210 16896 16526 16897
rect 16210 16832 16216 16896
rect 16280 16832 16296 16896
rect 16360 16832 16376 16896
rect 16440 16832 16456 16896
rect 16520 16832 16526 16896
rect 16210 16831 16526 16832
rect 7210 16352 7526 16353
rect 7210 16288 7216 16352
rect 7280 16288 7296 16352
rect 7360 16288 7376 16352
rect 7440 16288 7456 16352
rect 7520 16288 7526 16352
rect 7210 16287 7526 16288
rect 13210 16352 13526 16353
rect 13210 16288 13216 16352
rect 13280 16288 13296 16352
rect 13360 16288 13376 16352
rect 13440 16288 13456 16352
rect 13520 16288 13526 16352
rect 13210 16287 13526 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 10210 15808 10526 15809
rect 10210 15744 10216 15808
rect 10280 15744 10296 15808
rect 10360 15744 10376 15808
rect 10440 15744 10456 15808
rect 10520 15744 10526 15808
rect 10210 15743 10526 15744
rect 16210 15808 16526 15809
rect 16210 15744 16216 15808
rect 16280 15744 16296 15808
rect 16360 15744 16376 15808
rect 16440 15744 16456 15808
rect 16520 15744 16526 15808
rect 16210 15743 16526 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 7210 15264 7526 15265
rect 7210 15200 7216 15264
rect 7280 15200 7296 15264
rect 7360 15200 7376 15264
rect 7440 15200 7456 15264
rect 7520 15200 7526 15264
rect 7210 15199 7526 15200
rect 13210 15264 13526 15265
rect 13210 15200 13216 15264
rect 13280 15200 13296 15264
rect 13360 15200 13376 15264
rect 13440 15200 13456 15264
rect 13520 15200 13526 15264
rect 13210 15199 13526 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 10210 14720 10526 14721
rect 10210 14656 10216 14720
rect 10280 14656 10296 14720
rect 10360 14656 10376 14720
rect 10440 14656 10456 14720
rect 10520 14656 10526 14720
rect 10210 14655 10526 14656
rect 16210 14720 16526 14721
rect 16210 14656 16216 14720
rect 16280 14656 16296 14720
rect 16360 14656 16376 14720
rect 16440 14656 16456 14720
rect 16520 14656 16526 14720
rect 16210 14655 16526 14656
rect 7210 14176 7526 14177
rect 7210 14112 7216 14176
rect 7280 14112 7296 14176
rect 7360 14112 7376 14176
rect 7440 14112 7456 14176
rect 7520 14112 7526 14176
rect 7210 14111 7526 14112
rect 13210 14176 13526 14177
rect 13210 14112 13216 14176
rect 13280 14112 13296 14176
rect 13360 14112 13376 14176
rect 13440 14112 13456 14176
rect 13520 14112 13526 14176
rect 13210 14111 13526 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 10210 13632 10526 13633
rect 10210 13568 10216 13632
rect 10280 13568 10296 13632
rect 10360 13568 10376 13632
rect 10440 13568 10456 13632
rect 10520 13568 10526 13632
rect 10210 13567 10526 13568
rect 16210 13632 16526 13633
rect 16210 13568 16216 13632
rect 16280 13568 16296 13632
rect 16360 13568 16376 13632
rect 16440 13568 16456 13632
rect 16520 13568 16526 13632
rect 16210 13567 16526 13568
rect 7210 13088 7526 13089
rect 7210 13024 7216 13088
rect 7280 13024 7296 13088
rect 7360 13024 7376 13088
rect 7440 13024 7456 13088
rect 7520 13024 7526 13088
rect 7210 13023 7526 13024
rect 13210 13088 13526 13089
rect 13210 13024 13216 13088
rect 13280 13024 13296 13088
rect 13360 13024 13376 13088
rect 13440 13024 13456 13088
rect 13520 13024 13526 13088
rect 13210 13023 13526 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 10210 12544 10526 12545
rect 10210 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10526 12544
rect 10210 12479 10526 12480
rect 16210 12544 16526 12545
rect 16210 12480 16216 12544
rect 16280 12480 16296 12544
rect 16360 12480 16376 12544
rect 16440 12480 16456 12544
rect 16520 12480 16526 12544
rect 16210 12479 16526 12480
rect 16113 12338 16179 12341
rect 17506 12338 18306 12368
rect 16113 12336 18306 12338
rect 16113 12280 16118 12336
rect 16174 12280 18306 12336
rect 16113 12278 18306 12280
rect 16113 12275 16179 12278
rect 17506 12248 18306 12278
rect 7210 12000 7526 12001
rect 7210 11936 7216 12000
rect 7280 11936 7296 12000
rect 7360 11936 7376 12000
rect 7440 11936 7456 12000
rect 7520 11936 7526 12000
rect 7210 11935 7526 11936
rect 13210 12000 13526 12001
rect 13210 11936 13216 12000
rect 13280 11936 13296 12000
rect 13360 11936 13376 12000
rect 13440 11936 13456 12000
rect 13520 11936 13526 12000
rect 13210 11935 13526 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 10210 11456 10526 11457
rect 10210 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10526 11456
rect 10210 11391 10526 11392
rect 16210 11456 16526 11457
rect 16210 11392 16216 11456
rect 16280 11392 16296 11456
rect 16360 11392 16376 11456
rect 16440 11392 16456 11456
rect 16520 11392 16526 11456
rect 16210 11391 16526 11392
rect 7210 10912 7526 10913
rect 7210 10848 7216 10912
rect 7280 10848 7296 10912
rect 7360 10848 7376 10912
rect 7440 10848 7456 10912
rect 7520 10848 7526 10912
rect 7210 10847 7526 10848
rect 13210 10912 13526 10913
rect 13210 10848 13216 10912
rect 13280 10848 13296 10912
rect 13360 10848 13376 10912
rect 13440 10848 13456 10912
rect 13520 10848 13526 10912
rect 13210 10847 13526 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 10210 10368 10526 10369
rect 10210 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10526 10368
rect 10210 10303 10526 10304
rect 16210 10368 16526 10369
rect 16210 10304 16216 10368
rect 16280 10304 16296 10368
rect 16360 10304 16376 10368
rect 16440 10304 16456 10368
rect 16520 10304 16526 10368
rect 16210 10303 16526 10304
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10208 800 10238
rect 933 10235 999 10238
rect 7210 9824 7526 9825
rect 7210 9760 7216 9824
rect 7280 9760 7296 9824
rect 7360 9760 7376 9824
rect 7440 9760 7456 9824
rect 7520 9760 7526 9824
rect 7210 9759 7526 9760
rect 13210 9824 13526 9825
rect 13210 9760 13216 9824
rect 13280 9760 13296 9824
rect 13360 9760 13376 9824
rect 13440 9760 13456 9824
rect 13520 9760 13526 9824
rect 13210 9759 13526 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 10210 9280 10526 9281
rect 10210 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10526 9280
rect 10210 9215 10526 9216
rect 16210 9280 16526 9281
rect 16210 9216 16216 9280
rect 16280 9216 16296 9280
rect 16360 9216 16376 9280
rect 16440 9216 16456 9280
rect 16520 9216 16526 9280
rect 16210 9215 16526 9216
rect 7210 8736 7526 8737
rect 7210 8672 7216 8736
rect 7280 8672 7296 8736
rect 7360 8672 7376 8736
rect 7440 8672 7456 8736
rect 7520 8672 7526 8736
rect 7210 8671 7526 8672
rect 13210 8736 13526 8737
rect 13210 8672 13216 8736
rect 13280 8672 13296 8736
rect 13360 8672 13376 8736
rect 13440 8672 13456 8736
rect 13520 8672 13526 8736
rect 13210 8671 13526 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 10210 8192 10526 8193
rect 10210 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10526 8192
rect 10210 8127 10526 8128
rect 16210 8192 16526 8193
rect 16210 8128 16216 8192
rect 16280 8128 16296 8192
rect 16360 8128 16376 8192
rect 16440 8128 16456 8192
rect 16520 8128 16526 8192
rect 16210 8127 16526 8128
rect 7210 7648 7526 7649
rect 7210 7584 7216 7648
rect 7280 7584 7296 7648
rect 7360 7584 7376 7648
rect 7440 7584 7456 7648
rect 7520 7584 7526 7648
rect 7210 7583 7526 7584
rect 13210 7648 13526 7649
rect 13210 7584 13216 7648
rect 13280 7584 13296 7648
rect 13360 7584 13376 7648
rect 13440 7584 13456 7648
rect 13520 7584 13526 7648
rect 13210 7583 13526 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 10210 7104 10526 7105
rect 10210 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10526 7104
rect 10210 7039 10526 7040
rect 16210 7104 16526 7105
rect 16210 7040 16216 7104
rect 16280 7040 16296 7104
rect 16360 7040 16376 7104
rect 16440 7040 16456 7104
rect 16520 7040 16526 7104
rect 16210 7039 16526 7040
rect 17125 6898 17191 6901
rect 17506 6898 18306 6928
rect 17125 6896 18306 6898
rect 17125 6840 17130 6896
rect 17186 6840 18306 6896
rect 17125 6838 18306 6840
rect 17125 6835 17191 6838
rect 17506 6808 18306 6838
rect 7210 6560 7526 6561
rect 7210 6496 7216 6560
rect 7280 6496 7296 6560
rect 7360 6496 7376 6560
rect 7440 6496 7456 6560
rect 7520 6496 7526 6560
rect 7210 6495 7526 6496
rect 13210 6560 13526 6561
rect 13210 6496 13216 6560
rect 13280 6496 13296 6560
rect 13360 6496 13376 6560
rect 13440 6496 13456 6560
rect 13520 6496 13526 6560
rect 13210 6495 13526 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 10210 6016 10526 6017
rect 10210 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10526 6016
rect 10210 5951 10526 5952
rect 16210 6016 16526 6017
rect 16210 5952 16216 6016
rect 16280 5952 16296 6016
rect 16360 5952 16376 6016
rect 16440 5952 16456 6016
rect 16520 5952 16526 6016
rect 16210 5951 16526 5952
rect 7210 5472 7526 5473
rect 7210 5408 7216 5472
rect 7280 5408 7296 5472
rect 7360 5408 7376 5472
rect 7440 5408 7456 5472
rect 7520 5408 7526 5472
rect 7210 5407 7526 5408
rect 13210 5472 13526 5473
rect 13210 5408 13216 5472
rect 13280 5408 13296 5472
rect 13360 5408 13376 5472
rect 13440 5408 13456 5472
rect 13520 5408 13526 5472
rect 13210 5407 13526 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 10210 4928 10526 4929
rect 10210 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10526 4928
rect 10210 4863 10526 4864
rect 16210 4928 16526 4929
rect 16210 4864 16216 4928
rect 16280 4864 16296 4928
rect 16360 4864 16376 4928
rect 16440 4864 16456 4928
rect 16520 4864 16526 4928
rect 16210 4863 16526 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 7210 4384 7526 4385
rect 7210 4320 7216 4384
rect 7280 4320 7296 4384
rect 7360 4320 7376 4384
rect 7440 4320 7456 4384
rect 7520 4320 7526 4384
rect 7210 4319 7526 4320
rect 13210 4384 13526 4385
rect 13210 4320 13216 4384
rect 13280 4320 13296 4384
rect 13360 4320 13376 4384
rect 13440 4320 13456 4384
rect 13520 4320 13526 4384
rect 13210 4319 13526 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 10210 3840 10526 3841
rect 10210 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10526 3840
rect 10210 3775 10526 3776
rect 16210 3840 16526 3841
rect 16210 3776 16216 3840
rect 16280 3776 16296 3840
rect 16360 3776 16376 3840
rect 16440 3776 16456 3840
rect 16520 3776 16526 3840
rect 16210 3775 16526 3776
rect 7210 3296 7526 3297
rect 7210 3232 7216 3296
rect 7280 3232 7296 3296
rect 7360 3232 7376 3296
rect 7440 3232 7456 3296
rect 7520 3232 7526 3296
rect 7210 3231 7526 3232
rect 13210 3296 13526 3297
rect 13210 3232 13216 3296
rect 13280 3232 13296 3296
rect 13360 3232 13376 3296
rect 13440 3232 13456 3296
rect 13520 3232 13526 3296
rect 13210 3231 13526 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 10210 2752 10526 2753
rect 10210 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10526 2752
rect 10210 2687 10526 2688
rect 16210 2752 16526 2753
rect 16210 2688 16216 2752
rect 16280 2688 16296 2752
rect 16360 2688 16376 2752
rect 16440 2688 16456 2752
rect 16520 2688 16526 2752
rect 16210 2687 16526 2688
rect 7210 2208 7526 2209
rect 7210 2144 7216 2208
rect 7280 2144 7296 2208
rect 7360 2144 7376 2208
rect 7440 2144 7456 2208
rect 7520 2144 7526 2208
rect 7210 2143 7526 2144
rect 13210 2208 13526 2209
rect 13210 2144 13216 2208
rect 13280 2144 13296 2208
rect 13360 2144 13376 2208
rect 13440 2144 13456 2208
rect 13520 2144 13526 2208
rect 13210 2143 13526 2144
rect 17033 1458 17099 1461
rect 17506 1458 18306 1488
rect 17033 1456 18306 1458
rect 17033 1400 17038 1456
rect 17094 1400 18306 1456
rect 17033 1398 18306 1400
rect 17033 1395 17099 1398
rect 17506 1368 18306 1398
<< via3 >>
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 10216 17980 10280 17984
rect 10216 17924 10220 17980
rect 10220 17924 10276 17980
rect 10276 17924 10280 17980
rect 10216 17920 10280 17924
rect 10296 17980 10360 17984
rect 10296 17924 10300 17980
rect 10300 17924 10356 17980
rect 10356 17924 10360 17980
rect 10296 17920 10360 17924
rect 10376 17980 10440 17984
rect 10376 17924 10380 17980
rect 10380 17924 10436 17980
rect 10436 17924 10440 17980
rect 10376 17920 10440 17924
rect 10456 17980 10520 17984
rect 10456 17924 10460 17980
rect 10460 17924 10516 17980
rect 10516 17924 10520 17980
rect 10456 17920 10520 17924
rect 16216 17980 16280 17984
rect 16216 17924 16220 17980
rect 16220 17924 16276 17980
rect 16276 17924 16280 17980
rect 16216 17920 16280 17924
rect 16296 17980 16360 17984
rect 16296 17924 16300 17980
rect 16300 17924 16356 17980
rect 16356 17924 16360 17980
rect 16296 17920 16360 17924
rect 16376 17980 16440 17984
rect 16376 17924 16380 17980
rect 16380 17924 16436 17980
rect 16436 17924 16440 17980
rect 16376 17920 16440 17924
rect 16456 17980 16520 17984
rect 16456 17924 16460 17980
rect 16460 17924 16516 17980
rect 16516 17924 16520 17980
rect 16456 17920 16520 17924
rect 7216 17436 7280 17440
rect 7216 17380 7220 17436
rect 7220 17380 7276 17436
rect 7276 17380 7280 17436
rect 7216 17376 7280 17380
rect 7296 17436 7360 17440
rect 7296 17380 7300 17436
rect 7300 17380 7356 17436
rect 7356 17380 7360 17436
rect 7296 17376 7360 17380
rect 7376 17436 7440 17440
rect 7376 17380 7380 17436
rect 7380 17380 7436 17436
rect 7436 17380 7440 17436
rect 7376 17376 7440 17380
rect 7456 17436 7520 17440
rect 7456 17380 7460 17436
rect 7460 17380 7516 17436
rect 7516 17380 7520 17436
rect 7456 17376 7520 17380
rect 13216 17436 13280 17440
rect 13216 17380 13220 17436
rect 13220 17380 13276 17436
rect 13276 17380 13280 17436
rect 13216 17376 13280 17380
rect 13296 17436 13360 17440
rect 13296 17380 13300 17436
rect 13300 17380 13356 17436
rect 13356 17380 13360 17436
rect 13296 17376 13360 17380
rect 13376 17436 13440 17440
rect 13376 17380 13380 17436
rect 13380 17380 13436 17436
rect 13436 17380 13440 17436
rect 13376 17376 13440 17380
rect 13456 17436 13520 17440
rect 13456 17380 13460 17436
rect 13460 17380 13516 17436
rect 13516 17380 13520 17436
rect 13456 17376 13520 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 10216 16892 10280 16896
rect 10216 16836 10220 16892
rect 10220 16836 10276 16892
rect 10276 16836 10280 16892
rect 10216 16832 10280 16836
rect 10296 16892 10360 16896
rect 10296 16836 10300 16892
rect 10300 16836 10356 16892
rect 10356 16836 10360 16892
rect 10296 16832 10360 16836
rect 10376 16892 10440 16896
rect 10376 16836 10380 16892
rect 10380 16836 10436 16892
rect 10436 16836 10440 16892
rect 10376 16832 10440 16836
rect 10456 16892 10520 16896
rect 10456 16836 10460 16892
rect 10460 16836 10516 16892
rect 10516 16836 10520 16892
rect 10456 16832 10520 16836
rect 16216 16892 16280 16896
rect 16216 16836 16220 16892
rect 16220 16836 16276 16892
rect 16276 16836 16280 16892
rect 16216 16832 16280 16836
rect 16296 16892 16360 16896
rect 16296 16836 16300 16892
rect 16300 16836 16356 16892
rect 16356 16836 16360 16892
rect 16296 16832 16360 16836
rect 16376 16892 16440 16896
rect 16376 16836 16380 16892
rect 16380 16836 16436 16892
rect 16436 16836 16440 16892
rect 16376 16832 16440 16836
rect 16456 16892 16520 16896
rect 16456 16836 16460 16892
rect 16460 16836 16516 16892
rect 16516 16836 16520 16892
rect 16456 16832 16520 16836
rect 7216 16348 7280 16352
rect 7216 16292 7220 16348
rect 7220 16292 7276 16348
rect 7276 16292 7280 16348
rect 7216 16288 7280 16292
rect 7296 16348 7360 16352
rect 7296 16292 7300 16348
rect 7300 16292 7356 16348
rect 7356 16292 7360 16348
rect 7296 16288 7360 16292
rect 7376 16348 7440 16352
rect 7376 16292 7380 16348
rect 7380 16292 7436 16348
rect 7436 16292 7440 16348
rect 7376 16288 7440 16292
rect 7456 16348 7520 16352
rect 7456 16292 7460 16348
rect 7460 16292 7516 16348
rect 7516 16292 7520 16348
rect 7456 16288 7520 16292
rect 13216 16348 13280 16352
rect 13216 16292 13220 16348
rect 13220 16292 13276 16348
rect 13276 16292 13280 16348
rect 13216 16288 13280 16292
rect 13296 16348 13360 16352
rect 13296 16292 13300 16348
rect 13300 16292 13356 16348
rect 13356 16292 13360 16348
rect 13296 16288 13360 16292
rect 13376 16348 13440 16352
rect 13376 16292 13380 16348
rect 13380 16292 13436 16348
rect 13436 16292 13440 16348
rect 13376 16288 13440 16292
rect 13456 16348 13520 16352
rect 13456 16292 13460 16348
rect 13460 16292 13516 16348
rect 13516 16292 13520 16348
rect 13456 16288 13520 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 10216 15804 10280 15808
rect 10216 15748 10220 15804
rect 10220 15748 10276 15804
rect 10276 15748 10280 15804
rect 10216 15744 10280 15748
rect 10296 15804 10360 15808
rect 10296 15748 10300 15804
rect 10300 15748 10356 15804
rect 10356 15748 10360 15804
rect 10296 15744 10360 15748
rect 10376 15804 10440 15808
rect 10376 15748 10380 15804
rect 10380 15748 10436 15804
rect 10436 15748 10440 15804
rect 10376 15744 10440 15748
rect 10456 15804 10520 15808
rect 10456 15748 10460 15804
rect 10460 15748 10516 15804
rect 10516 15748 10520 15804
rect 10456 15744 10520 15748
rect 16216 15804 16280 15808
rect 16216 15748 16220 15804
rect 16220 15748 16276 15804
rect 16276 15748 16280 15804
rect 16216 15744 16280 15748
rect 16296 15804 16360 15808
rect 16296 15748 16300 15804
rect 16300 15748 16356 15804
rect 16356 15748 16360 15804
rect 16296 15744 16360 15748
rect 16376 15804 16440 15808
rect 16376 15748 16380 15804
rect 16380 15748 16436 15804
rect 16436 15748 16440 15804
rect 16376 15744 16440 15748
rect 16456 15804 16520 15808
rect 16456 15748 16460 15804
rect 16460 15748 16516 15804
rect 16516 15748 16520 15804
rect 16456 15744 16520 15748
rect 7216 15260 7280 15264
rect 7216 15204 7220 15260
rect 7220 15204 7276 15260
rect 7276 15204 7280 15260
rect 7216 15200 7280 15204
rect 7296 15260 7360 15264
rect 7296 15204 7300 15260
rect 7300 15204 7356 15260
rect 7356 15204 7360 15260
rect 7296 15200 7360 15204
rect 7376 15260 7440 15264
rect 7376 15204 7380 15260
rect 7380 15204 7436 15260
rect 7436 15204 7440 15260
rect 7376 15200 7440 15204
rect 7456 15260 7520 15264
rect 7456 15204 7460 15260
rect 7460 15204 7516 15260
rect 7516 15204 7520 15260
rect 7456 15200 7520 15204
rect 13216 15260 13280 15264
rect 13216 15204 13220 15260
rect 13220 15204 13276 15260
rect 13276 15204 13280 15260
rect 13216 15200 13280 15204
rect 13296 15260 13360 15264
rect 13296 15204 13300 15260
rect 13300 15204 13356 15260
rect 13356 15204 13360 15260
rect 13296 15200 13360 15204
rect 13376 15260 13440 15264
rect 13376 15204 13380 15260
rect 13380 15204 13436 15260
rect 13436 15204 13440 15260
rect 13376 15200 13440 15204
rect 13456 15260 13520 15264
rect 13456 15204 13460 15260
rect 13460 15204 13516 15260
rect 13516 15204 13520 15260
rect 13456 15200 13520 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 10216 14716 10280 14720
rect 10216 14660 10220 14716
rect 10220 14660 10276 14716
rect 10276 14660 10280 14716
rect 10216 14656 10280 14660
rect 10296 14716 10360 14720
rect 10296 14660 10300 14716
rect 10300 14660 10356 14716
rect 10356 14660 10360 14716
rect 10296 14656 10360 14660
rect 10376 14716 10440 14720
rect 10376 14660 10380 14716
rect 10380 14660 10436 14716
rect 10436 14660 10440 14716
rect 10376 14656 10440 14660
rect 10456 14716 10520 14720
rect 10456 14660 10460 14716
rect 10460 14660 10516 14716
rect 10516 14660 10520 14716
rect 10456 14656 10520 14660
rect 16216 14716 16280 14720
rect 16216 14660 16220 14716
rect 16220 14660 16276 14716
rect 16276 14660 16280 14716
rect 16216 14656 16280 14660
rect 16296 14716 16360 14720
rect 16296 14660 16300 14716
rect 16300 14660 16356 14716
rect 16356 14660 16360 14716
rect 16296 14656 16360 14660
rect 16376 14716 16440 14720
rect 16376 14660 16380 14716
rect 16380 14660 16436 14716
rect 16436 14660 16440 14716
rect 16376 14656 16440 14660
rect 16456 14716 16520 14720
rect 16456 14660 16460 14716
rect 16460 14660 16516 14716
rect 16516 14660 16520 14716
rect 16456 14656 16520 14660
rect 7216 14172 7280 14176
rect 7216 14116 7220 14172
rect 7220 14116 7276 14172
rect 7276 14116 7280 14172
rect 7216 14112 7280 14116
rect 7296 14172 7360 14176
rect 7296 14116 7300 14172
rect 7300 14116 7356 14172
rect 7356 14116 7360 14172
rect 7296 14112 7360 14116
rect 7376 14172 7440 14176
rect 7376 14116 7380 14172
rect 7380 14116 7436 14172
rect 7436 14116 7440 14172
rect 7376 14112 7440 14116
rect 7456 14172 7520 14176
rect 7456 14116 7460 14172
rect 7460 14116 7516 14172
rect 7516 14116 7520 14172
rect 7456 14112 7520 14116
rect 13216 14172 13280 14176
rect 13216 14116 13220 14172
rect 13220 14116 13276 14172
rect 13276 14116 13280 14172
rect 13216 14112 13280 14116
rect 13296 14172 13360 14176
rect 13296 14116 13300 14172
rect 13300 14116 13356 14172
rect 13356 14116 13360 14172
rect 13296 14112 13360 14116
rect 13376 14172 13440 14176
rect 13376 14116 13380 14172
rect 13380 14116 13436 14172
rect 13436 14116 13440 14172
rect 13376 14112 13440 14116
rect 13456 14172 13520 14176
rect 13456 14116 13460 14172
rect 13460 14116 13516 14172
rect 13516 14116 13520 14172
rect 13456 14112 13520 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 10216 13628 10280 13632
rect 10216 13572 10220 13628
rect 10220 13572 10276 13628
rect 10276 13572 10280 13628
rect 10216 13568 10280 13572
rect 10296 13628 10360 13632
rect 10296 13572 10300 13628
rect 10300 13572 10356 13628
rect 10356 13572 10360 13628
rect 10296 13568 10360 13572
rect 10376 13628 10440 13632
rect 10376 13572 10380 13628
rect 10380 13572 10436 13628
rect 10436 13572 10440 13628
rect 10376 13568 10440 13572
rect 10456 13628 10520 13632
rect 10456 13572 10460 13628
rect 10460 13572 10516 13628
rect 10516 13572 10520 13628
rect 10456 13568 10520 13572
rect 16216 13628 16280 13632
rect 16216 13572 16220 13628
rect 16220 13572 16276 13628
rect 16276 13572 16280 13628
rect 16216 13568 16280 13572
rect 16296 13628 16360 13632
rect 16296 13572 16300 13628
rect 16300 13572 16356 13628
rect 16356 13572 16360 13628
rect 16296 13568 16360 13572
rect 16376 13628 16440 13632
rect 16376 13572 16380 13628
rect 16380 13572 16436 13628
rect 16436 13572 16440 13628
rect 16376 13568 16440 13572
rect 16456 13628 16520 13632
rect 16456 13572 16460 13628
rect 16460 13572 16516 13628
rect 16516 13572 16520 13628
rect 16456 13568 16520 13572
rect 7216 13084 7280 13088
rect 7216 13028 7220 13084
rect 7220 13028 7276 13084
rect 7276 13028 7280 13084
rect 7216 13024 7280 13028
rect 7296 13084 7360 13088
rect 7296 13028 7300 13084
rect 7300 13028 7356 13084
rect 7356 13028 7360 13084
rect 7296 13024 7360 13028
rect 7376 13084 7440 13088
rect 7376 13028 7380 13084
rect 7380 13028 7436 13084
rect 7436 13028 7440 13084
rect 7376 13024 7440 13028
rect 7456 13084 7520 13088
rect 7456 13028 7460 13084
rect 7460 13028 7516 13084
rect 7516 13028 7520 13084
rect 7456 13024 7520 13028
rect 13216 13084 13280 13088
rect 13216 13028 13220 13084
rect 13220 13028 13276 13084
rect 13276 13028 13280 13084
rect 13216 13024 13280 13028
rect 13296 13084 13360 13088
rect 13296 13028 13300 13084
rect 13300 13028 13356 13084
rect 13356 13028 13360 13084
rect 13296 13024 13360 13028
rect 13376 13084 13440 13088
rect 13376 13028 13380 13084
rect 13380 13028 13436 13084
rect 13436 13028 13440 13084
rect 13376 13024 13440 13028
rect 13456 13084 13520 13088
rect 13456 13028 13460 13084
rect 13460 13028 13516 13084
rect 13516 13028 13520 13084
rect 13456 13024 13520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 10216 12540 10280 12544
rect 10216 12484 10220 12540
rect 10220 12484 10276 12540
rect 10276 12484 10280 12540
rect 10216 12480 10280 12484
rect 10296 12540 10360 12544
rect 10296 12484 10300 12540
rect 10300 12484 10356 12540
rect 10356 12484 10360 12540
rect 10296 12480 10360 12484
rect 10376 12540 10440 12544
rect 10376 12484 10380 12540
rect 10380 12484 10436 12540
rect 10436 12484 10440 12540
rect 10376 12480 10440 12484
rect 10456 12540 10520 12544
rect 10456 12484 10460 12540
rect 10460 12484 10516 12540
rect 10516 12484 10520 12540
rect 10456 12480 10520 12484
rect 16216 12540 16280 12544
rect 16216 12484 16220 12540
rect 16220 12484 16276 12540
rect 16276 12484 16280 12540
rect 16216 12480 16280 12484
rect 16296 12540 16360 12544
rect 16296 12484 16300 12540
rect 16300 12484 16356 12540
rect 16356 12484 16360 12540
rect 16296 12480 16360 12484
rect 16376 12540 16440 12544
rect 16376 12484 16380 12540
rect 16380 12484 16436 12540
rect 16436 12484 16440 12540
rect 16376 12480 16440 12484
rect 16456 12540 16520 12544
rect 16456 12484 16460 12540
rect 16460 12484 16516 12540
rect 16516 12484 16520 12540
rect 16456 12480 16520 12484
rect 7216 11996 7280 12000
rect 7216 11940 7220 11996
rect 7220 11940 7276 11996
rect 7276 11940 7280 11996
rect 7216 11936 7280 11940
rect 7296 11996 7360 12000
rect 7296 11940 7300 11996
rect 7300 11940 7356 11996
rect 7356 11940 7360 11996
rect 7296 11936 7360 11940
rect 7376 11996 7440 12000
rect 7376 11940 7380 11996
rect 7380 11940 7436 11996
rect 7436 11940 7440 11996
rect 7376 11936 7440 11940
rect 7456 11996 7520 12000
rect 7456 11940 7460 11996
rect 7460 11940 7516 11996
rect 7516 11940 7520 11996
rect 7456 11936 7520 11940
rect 13216 11996 13280 12000
rect 13216 11940 13220 11996
rect 13220 11940 13276 11996
rect 13276 11940 13280 11996
rect 13216 11936 13280 11940
rect 13296 11996 13360 12000
rect 13296 11940 13300 11996
rect 13300 11940 13356 11996
rect 13356 11940 13360 11996
rect 13296 11936 13360 11940
rect 13376 11996 13440 12000
rect 13376 11940 13380 11996
rect 13380 11940 13436 11996
rect 13436 11940 13440 11996
rect 13376 11936 13440 11940
rect 13456 11996 13520 12000
rect 13456 11940 13460 11996
rect 13460 11940 13516 11996
rect 13516 11940 13520 11996
rect 13456 11936 13520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 10216 11452 10280 11456
rect 10216 11396 10220 11452
rect 10220 11396 10276 11452
rect 10276 11396 10280 11452
rect 10216 11392 10280 11396
rect 10296 11452 10360 11456
rect 10296 11396 10300 11452
rect 10300 11396 10356 11452
rect 10356 11396 10360 11452
rect 10296 11392 10360 11396
rect 10376 11452 10440 11456
rect 10376 11396 10380 11452
rect 10380 11396 10436 11452
rect 10436 11396 10440 11452
rect 10376 11392 10440 11396
rect 10456 11452 10520 11456
rect 10456 11396 10460 11452
rect 10460 11396 10516 11452
rect 10516 11396 10520 11452
rect 10456 11392 10520 11396
rect 16216 11452 16280 11456
rect 16216 11396 16220 11452
rect 16220 11396 16276 11452
rect 16276 11396 16280 11452
rect 16216 11392 16280 11396
rect 16296 11452 16360 11456
rect 16296 11396 16300 11452
rect 16300 11396 16356 11452
rect 16356 11396 16360 11452
rect 16296 11392 16360 11396
rect 16376 11452 16440 11456
rect 16376 11396 16380 11452
rect 16380 11396 16436 11452
rect 16436 11396 16440 11452
rect 16376 11392 16440 11396
rect 16456 11452 16520 11456
rect 16456 11396 16460 11452
rect 16460 11396 16516 11452
rect 16516 11396 16520 11452
rect 16456 11392 16520 11396
rect 7216 10908 7280 10912
rect 7216 10852 7220 10908
rect 7220 10852 7276 10908
rect 7276 10852 7280 10908
rect 7216 10848 7280 10852
rect 7296 10908 7360 10912
rect 7296 10852 7300 10908
rect 7300 10852 7356 10908
rect 7356 10852 7360 10908
rect 7296 10848 7360 10852
rect 7376 10908 7440 10912
rect 7376 10852 7380 10908
rect 7380 10852 7436 10908
rect 7436 10852 7440 10908
rect 7376 10848 7440 10852
rect 7456 10908 7520 10912
rect 7456 10852 7460 10908
rect 7460 10852 7516 10908
rect 7516 10852 7520 10908
rect 7456 10848 7520 10852
rect 13216 10908 13280 10912
rect 13216 10852 13220 10908
rect 13220 10852 13276 10908
rect 13276 10852 13280 10908
rect 13216 10848 13280 10852
rect 13296 10908 13360 10912
rect 13296 10852 13300 10908
rect 13300 10852 13356 10908
rect 13356 10852 13360 10908
rect 13296 10848 13360 10852
rect 13376 10908 13440 10912
rect 13376 10852 13380 10908
rect 13380 10852 13436 10908
rect 13436 10852 13440 10908
rect 13376 10848 13440 10852
rect 13456 10908 13520 10912
rect 13456 10852 13460 10908
rect 13460 10852 13516 10908
rect 13516 10852 13520 10908
rect 13456 10848 13520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 10216 10364 10280 10368
rect 10216 10308 10220 10364
rect 10220 10308 10276 10364
rect 10276 10308 10280 10364
rect 10216 10304 10280 10308
rect 10296 10364 10360 10368
rect 10296 10308 10300 10364
rect 10300 10308 10356 10364
rect 10356 10308 10360 10364
rect 10296 10304 10360 10308
rect 10376 10364 10440 10368
rect 10376 10308 10380 10364
rect 10380 10308 10436 10364
rect 10436 10308 10440 10364
rect 10376 10304 10440 10308
rect 10456 10364 10520 10368
rect 10456 10308 10460 10364
rect 10460 10308 10516 10364
rect 10516 10308 10520 10364
rect 10456 10304 10520 10308
rect 16216 10364 16280 10368
rect 16216 10308 16220 10364
rect 16220 10308 16276 10364
rect 16276 10308 16280 10364
rect 16216 10304 16280 10308
rect 16296 10364 16360 10368
rect 16296 10308 16300 10364
rect 16300 10308 16356 10364
rect 16356 10308 16360 10364
rect 16296 10304 16360 10308
rect 16376 10364 16440 10368
rect 16376 10308 16380 10364
rect 16380 10308 16436 10364
rect 16436 10308 16440 10364
rect 16376 10304 16440 10308
rect 16456 10364 16520 10368
rect 16456 10308 16460 10364
rect 16460 10308 16516 10364
rect 16516 10308 16520 10364
rect 16456 10304 16520 10308
rect 7216 9820 7280 9824
rect 7216 9764 7220 9820
rect 7220 9764 7276 9820
rect 7276 9764 7280 9820
rect 7216 9760 7280 9764
rect 7296 9820 7360 9824
rect 7296 9764 7300 9820
rect 7300 9764 7356 9820
rect 7356 9764 7360 9820
rect 7296 9760 7360 9764
rect 7376 9820 7440 9824
rect 7376 9764 7380 9820
rect 7380 9764 7436 9820
rect 7436 9764 7440 9820
rect 7376 9760 7440 9764
rect 7456 9820 7520 9824
rect 7456 9764 7460 9820
rect 7460 9764 7516 9820
rect 7516 9764 7520 9820
rect 7456 9760 7520 9764
rect 13216 9820 13280 9824
rect 13216 9764 13220 9820
rect 13220 9764 13276 9820
rect 13276 9764 13280 9820
rect 13216 9760 13280 9764
rect 13296 9820 13360 9824
rect 13296 9764 13300 9820
rect 13300 9764 13356 9820
rect 13356 9764 13360 9820
rect 13296 9760 13360 9764
rect 13376 9820 13440 9824
rect 13376 9764 13380 9820
rect 13380 9764 13436 9820
rect 13436 9764 13440 9820
rect 13376 9760 13440 9764
rect 13456 9820 13520 9824
rect 13456 9764 13460 9820
rect 13460 9764 13516 9820
rect 13516 9764 13520 9820
rect 13456 9760 13520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 10216 9276 10280 9280
rect 10216 9220 10220 9276
rect 10220 9220 10276 9276
rect 10276 9220 10280 9276
rect 10216 9216 10280 9220
rect 10296 9276 10360 9280
rect 10296 9220 10300 9276
rect 10300 9220 10356 9276
rect 10356 9220 10360 9276
rect 10296 9216 10360 9220
rect 10376 9276 10440 9280
rect 10376 9220 10380 9276
rect 10380 9220 10436 9276
rect 10436 9220 10440 9276
rect 10376 9216 10440 9220
rect 10456 9276 10520 9280
rect 10456 9220 10460 9276
rect 10460 9220 10516 9276
rect 10516 9220 10520 9276
rect 10456 9216 10520 9220
rect 16216 9276 16280 9280
rect 16216 9220 16220 9276
rect 16220 9220 16276 9276
rect 16276 9220 16280 9276
rect 16216 9216 16280 9220
rect 16296 9276 16360 9280
rect 16296 9220 16300 9276
rect 16300 9220 16356 9276
rect 16356 9220 16360 9276
rect 16296 9216 16360 9220
rect 16376 9276 16440 9280
rect 16376 9220 16380 9276
rect 16380 9220 16436 9276
rect 16436 9220 16440 9276
rect 16376 9216 16440 9220
rect 16456 9276 16520 9280
rect 16456 9220 16460 9276
rect 16460 9220 16516 9276
rect 16516 9220 16520 9276
rect 16456 9216 16520 9220
rect 7216 8732 7280 8736
rect 7216 8676 7220 8732
rect 7220 8676 7276 8732
rect 7276 8676 7280 8732
rect 7216 8672 7280 8676
rect 7296 8732 7360 8736
rect 7296 8676 7300 8732
rect 7300 8676 7356 8732
rect 7356 8676 7360 8732
rect 7296 8672 7360 8676
rect 7376 8732 7440 8736
rect 7376 8676 7380 8732
rect 7380 8676 7436 8732
rect 7436 8676 7440 8732
rect 7376 8672 7440 8676
rect 7456 8732 7520 8736
rect 7456 8676 7460 8732
rect 7460 8676 7516 8732
rect 7516 8676 7520 8732
rect 7456 8672 7520 8676
rect 13216 8732 13280 8736
rect 13216 8676 13220 8732
rect 13220 8676 13276 8732
rect 13276 8676 13280 8732
rect 13216 8672 13280 8676
rect 13296 8732 13360 8736
rect 13296 8676 13300 8732
rect 13300 8676 13356 8732
rect 13356 8676 13360 8732
rect 13296 8672 13360 8676
rect 13376 8732 13440 8736
rect 13376 8676 13380 8732
rect 13380 8676 13436 8732
rect 13436 8676 13440 8732
rect 13376 8672 13440 8676
rect 13456 8732 13520 8736
rect 13456 8676 13460 8732
rect 13460 8676 13516 8732
rect 13516 8676 13520 8732
rect 13456 8672 13520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 10216 8188 10280 8192
rect 10216 8132 10220 8188
rect 10220 8132 10276 8188
rect 10276 8132 10280 8188
rect 10216 8128 10280 8132
rect 10296 8188 10360 8192
rect 10296 8132 10300 8188
rect 10300 8132 10356 8188
rect 10356 8132 10360 8188
rect 10296 8128 10360 8132
rect 10376 8188 10440 8192
rect 10376 8132 10380 8188
rect 10380 8132 10436 8188
rect 10436 8132 10440 8188
rect 10376 8128 10440 8132
rect 10456 8188 10520 8192
rect 10456 8132 10460 8188
rect 10460 8132 10516 8188
rect 10516 8132 10520 8188
rect 10456 8128 10520 8132
rect 16216 8188 16280 8192
rect 16216 8132 16220 8188
rect 16220 8132 16276 8188
rect 16276 8132 16280 8188
rect 16216 8128 16280 8132
rect 16296 8188 16360 8192
rect 16296 8132 16300 8188
rect 16300 8132 16356 8188
rect 16356 8132 16360 8188
rect 16296 8128 16360 8132
rect 16376 8188 16440 8192
rect 16376 8132 16380 8188
rect 16380 8132 16436 8188
rect 16436 8132 16440 8188
rect 16376 8128 16440 8132
rect 16456 8188 16520 8192
rect 16456 8132 16460 8188
rect 16460 8132 16516 8188
rect 16516 8132 16520 8188
rect 16456 8128 16520 8132
rect 7216 7644 7280 7648
rect 7216 7588 7220 7644
rect 7220 7588 7276 7644
rect 7276 7588 7280 7644
rect 7216 7584 7280 7588
rect 7296 7644 7360 7648
rect 7296 7588 7300 7644
rect 7300 7588 7356 7644
rect 7356 7588 7360 7644
rect 7296 7584 7360 7588
rect 7376 7644 7440 7648
rect 7376 7588 7380 7644
rect 7380 7588 7436 7644
rect 7436 7588 7440 7644
rect 7376 7584 7440 7588
rect 7456 7644 7520 7648
rect 7456 7588 7460 7644
rect 7460 7588 7516 7644
rect 7516 7588 7520 7644
rect 7456 7584 7520 7588
rect 13216 7644 13280 7648
rect 13216 7588 13220 7644
rect 13220 7588 13276 7644
rect 13276 7588 13280 7644
rect 13216 7584 13280 7588
rect 13296 7644 13360 7648
rect 13296 7588 13300 7644
rect 13300 7588 13356 7644
rect 13356 7588 13360 7644
rect 13296 7584 13360 7588
rect 13376 7644 13440 7648
rect 13376 7588 13380 7644
rect 13380 7588 13436 7644
rect 13436 7588 13440 7644
rect 13376 7584 13440 7588
rect 13456 7644 13520 7648
rect 13456 7588 13460 7644
rect 13460 7588 13516 7644
rect 13516 7588 13520 7644
rect 13456 7584 13520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 10216 7100 10280 7104
rect 10216 7044 10220 7100
rect 10220 7044 10276 7100
rect 10276 7044 10280 7100
rect 10216 7040 10280 7044
rect 10296 7100 10360 7104
rect 10296 7044 10300 7100
rect 10300 7044 10356 7100
rect 10356 7044 10360 7100
rect 10296 7040 10360 7044
rect 10376 7100 10440 7104
rect 10376 7044 10380 7100
rect 10380 7044 10436 7100
rect 10436 7044 10440 7100
rect 10376 7040 10440 7044
rect 10456 7100 10520 7104
rect 10456 7044 10460 7100
rect 10460 7044 10516 7100
rect 10516 7044 10520 7100
rect 10456 7040 10520 7044
rect 16216 7100 16280 7104
rect 16216 7044 16220 7100
rect 16220 7044 16276 7100
rect 16276 7044 16280 7100
rect 16216 7040 16280 7044
rect 16296 7100 16360 7104
rect 16296 7044 16300 7100
rect 16300 7044 16356 7100
rect 16356 7044 16360 7100
rect 16296 7040 16360 7044
rect 16376 7100 16440 7104
rect 16376 7044 16380 7100
rect 16380 7044 16436 7100
rect 16436 7044 16440 7100
rect 16376 7040 16440 7044
rect 16456 7100 16520 7104
rect 16456 7044 16460 7100
rect 16460 7044 16516 7100
rect 16516 7044 16520 7100
rect 16456 7040 16520 7044
rect 7216 6556 7280 6560
rect 7216 6500 7220 6556
rect 7220 6500 7276 6556
rect 7276 6500 7280 6556
rect 7216 6496 7280 6500
rect 7296 6556 7360 6560
rect 7296 6500 7300 6556
rect 7300 6500 7356 6556
rect 7356 6500 7360 6556
rect 7296 6496 7360 6500
rect 7376 6556 7440 6560
rect 7376 6500 7380 6556
rect 7380 6500 7436 6556
rect 7436 6500 7440 6556
rect 7376 6496 7440 6500
rect 7456 6556 7520 6560
rect 7456 6500 7460 6556
rect 7460 6500 7516 6556
rect 7516 6500 7520 6556
rect 7456 6496 7520 6500
rect 13216 6556 13280 6560
rect 13216 6500 13220 6556
rect 13220 6500 13276 6556
rect 13276 6500 13280 6556
rect 13216 6496 13280 6500
rect 13296 6556 13360 6560
rect 13296 6500 13300 6556
rect 13300 6500 13356 6556
rect 13356 6500 13360 6556
rect 13296 6496 13360 6500
rect 13376 6556 13440 6560
rect 13376 6500 13380 6556
rect 13380 6500 13436 6556
rect 13436 6500 13440 6556
rect 13376 6496 13440 6500
rect 13456 6556 13520 6560
rect 13456 6500 13460 6556
rect 13460 6500 13516 6556
rect 13516 6500 13520 6556
rect 13456 6496 13520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 10216 6012 10280 6016
rect 10216 5956 10220 6012
rect 10220 5956 10276 6012
rect 10276 5956 10280 6012
rect 10216 5952 10280 5956
rect 10296 6012 10360 6016
rect 10296 5956 10300 6012
rect 10300 5956 10356 6012
rect 10356 5956 10360 6012
rect 10296 5952 10360 5956
rect 10376 6012 10440 6016
rect 10376 5956 10380 6012
rect 10380 5956 10436 6012
rect 10436 5956 10440 6012
rect 10376 5952 10440 5956
rect 10456 6012 10520 6016
rect 10456 5956 10460 6012
rect 10460 5956 10516 6012
rect 10516 5956 10520 6012
rect 10456 5952 10520 5956
rect 16216 6012 16280 6016
rect 16216 5956 16220 6012
rect 16220 5956 16276 6012
rect 16276 5956 16280 6012
rect 16216 5952 16280 5956
rect 16296 6012 16360 6016
rect 16296 5956 16300 6012
rect 16300 5956 16356 6012
rect 16356 5956 16360 6012
rect 16296 5952 16360 5956
rect 16376 6012 16440 6016
rect 16376 5956 16380 6012
rect 16380 5956 16436 6012
rect 16436 5956 16440 6012
rect 16376 5952 16440 5956
rect 16456 6012 16520 6016
rect 16456 5956 16460 6012
rect 16460 5956 16516 6012
rect 16516 5956 16520 6012
rect 16456 5952 16520 5956
rect 7216 5468 7280 5472
rect 7216 5412 7220 5468
rect 7220 5412 7276 5468
rect 7276 5412 7280 5468
rect 7216 5408 7280 5412
rect 7296 5468 7360 5472
rect 7296 5412 7300 5468
rect 7300 5412 7356 5468
rect 7356 5412 7360 5468
rect 7296 5408 7360 5412
rect 7376 5468 7440 5472
rect 7376 5412 7380 5468
rect 7380 5412 7436 5468
rect 7436 5412 7440 5468
rect 7376 5408 7440 5412
rect 7456 5468 7520 5472
rect 7456 5412 7460 5468
rect 7460 5412 7516 5468
rect 7516 5412 7520 5468
rect 7456 5408 7520 5412
rect 13216 5468 13280 5472
rect 13216 5412 13220 5468
rect 13220 5412 13276 5468
rect 13276 5412 13280 5468
rect 13216 5408 13280 5412
rect 13296 5468 13360 5472
rect 13296 5412 13300 5468
rect 13300 5412 13356 5468
rect 13356 5412 13360 5468
rect 13296 5408 13360 5412
rect 13376 5468 13440 5472
rect 13376 5412 13380 5468
rect 13380 5412 13436 5468
rect 13436 5412 13440 5468
rect 13376 5408 13440 5412
rect 13456 5468 13520 5472
rect 13456 5412 13460 5468
rect 13460 5412 13516 5468
rect 13516 5412 13520 5468
rect 13456 5408 13520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 10216 4924 10280 4928
rect 10216 4868 10220 4924
rect 10220 4868 10276 4924
rect 10276 4868 10280 4924
rect 10216 4864 10280 4868
rect 10296 4924 10360 4928
rect 10296 4868 10300 4924
rect 10300 4868 10356 4924
rect 10356 4868 10360 4924
rect 10296 4864 10360 4868
rect 10376 4924 10440 4928
rect 10376 4868 10380 4924
rect 10380 4868 10436 4924
rect 10436 4868 10440 4924
rect 10376 4864 10440 4868
rect 10456 4924 10520 4928
rect 10456 4868 10460 4924
rect 10460 4868 10516 4924
rect 10516 4868 10520 4924
rect 10456 4864 10520 4868
rect 16216 4924 16280 4928
rect 16216 4868 16220 4924
rect 16220 4868 16276 4924
rect 16276 4868 16280 4924
rect 16216 4864 16280 4868
rect 16296 4924 16360 4928
rect 16296 4868 16300 4924
rect 16300 4868 16356 4924
rect 16356 4868 16360 4924
rect 16296 4864 16360 4868
rect 16376 4924 16440 4928
rect 16376 4868 16380 4924
rect 16380 4868 16436 4924
rect 16436 4868 16440 4924
rect 16376 4864 16440 4868
rect 16456 4924 16520 4928
rect 16456 4868 16460 4924
rect 16460 4868 16516 4924
rect 16516 4868 16520 4924
rect 16456 4864 16520 4868
rect 7216 4380 7280 4384
rect 7216 4324 7220 4380
rect 7220 4324 7276 4380
rect 7276 4324 7280 4380
rect 7216 4320 7280 4324
rect 7296 4380 7360 4384
rect 7296 4324 7300 4380
rect 7300 4324 7356 4380
rect 7356 4324 7360 4380
rect 7296 4320 7360 4324
rect 7376 4380 7440 4384
rect 7376 4324 7380 4380
rect 7380 4324 7436 4380
rect 7436 4324 7440 4380
rect 7376 4320 7440 4324
rect 7456 4380 7520 4384
rect 7456 4324 7460 4380
rect 7460 4324 7516 4380
rect 7516 4324 7520 4380
rect 7456 4320 7520 4324
rect 13216 4380 13280 4384
rect 13216 4324 13220 4380
rect 13220 4324 13276 4380
rect 13276 4324 13280 4380
rect 13216 4320 13280 4324
rect 13296 4380 13360 4384
rect 13296 4324 13300 4380
rect 13300 4324 13356 4380
rect 13356 4324 13360 4380
rect 13296 4320 13360 4324
rect 13376 4380 13440 4384
rect 13376 4324 13380 4380
rect 13380 4324 13436 4380
rect 13436 4324 13440 4380
rect 13376 4320 13440 4324
rect 13456 4380 13520 4384
rect 13456 4324 13460 4380
rect 13460 4324 13516 4380
rect 13516 4324 13520 4380
rect 13456 4320 13520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 10216 3836 10280 3840
rect 10216 3780 10220 3836
rect 10220 3780 10276 3836
rect 10276 3780 10280 3836
rect 10216 3776 10280 3780
rect 10296 3836 10360 3840
rect 10296 3780 10300 3836
rect 10300 3780 10356 3836
rect 10356 3780 10360 3836
rect 10296 3776 10360 3780
rect 10376 3836 10440 3840
rect 10376 3780 10380 3836
rect 10380 3780 10436 3836
rect 10436 3780 10440 3836
rect 10376 3776 10440 3780
rect 10456 3836 10520 3840
rect 10456 3780 10460 3836
rect 10460 3780 10516 3836
rect 10516 3780 10520 3836
rect 10456 3776 10520 3780
rect 16216 3836 16280 3840
rect 16216 3780 16220 3836
rect 16220 3780 16276 3836
rect 16276 3780 16280 3836
rect 16216 3776 16280 3780
rect 16296 3836 16360 3840
rect 16296 3780 16300 3836
rect 16300 3780 16356 3836
rect 16356 3780 16360 3836
rect 16296 3776 16360 3780
rect 16376 3836 16440 3840
rect 16376 3780 16380 3836
rect 16380 3780 16436 3836
rect 16436 3780 16440 3836
rect 16376 3776 16440 3780
rect 16456 3836 16520 3840
rect 16456 3780 16460 3836
rect 16460 3780 16516 3836
rect 16516 3780 16520 3836
rect 16456 3776 16520 3780
rect 7216 3292 7280 3296
rect 7216 3236 7220 3292
rect 7220 3236 7276 3292
rect 7276 3236 7280 3292
rect 7216 3232 7280 3236
rect 7296 3292 7360 3296
rect 7296 3236 7300 3292
rect 7300 3236 7356 3292
rect 7356 3236 7360 3292
rect 7296 3232 7360 3236
rect 7376 3292 7440 3296
rect 7376 3236 7380 3292
rect 7380 3236 7436 3292
rect 7436 3236 7440 3292
rect 7376 3232 7440 3236
rect 7456 3292 7520 3296
rect 7456 3236 7460 3292
rect 7460 3236 7516 3292
rect 7516 3236 7520 3292
rect 7456 3232 7520 3236
rect 13216 3292 13280 3296
rect 13216 3236 13220 3292
rect 13220 3236 13276 3292
rect 13276 3236 13280 3292
rect 13216 3232 13280 3236
rect 13296 3292 13360 3296
rect 13296 3236 13300 3292
rect 13300 3236 13356 3292
rect 13356 3236 13360 3292
rect 13296 3232 13360 3236
rect 13376 3292 13440 3296
rect 13376 3236 13380 3292
rect 13380 3236 13436 3292
rect 13436 3236 13440 3292
rect 13376 3232 13440 3236
rect 13456 3292 13520 3296
rect 13456 3236 13460 3292
rect 13460 3236 13516 3292
rect 13516 3236 13520 3292
rect 13456 3232 13520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 10216 2748 10280 2752
rect 10216 2692 10220 2748
rect 10220 2692 10276 2748
rect 10276 2692 10280 2748
rect 10216 2688 10280 2692
rect 10296 2748 10360 2752
rect 10296 2692 10300 2748
rect 10300 2692 10356 2748
rect 10356 2692 10360 2748
rect 10296 2688 10360 2692
rect 10376 2748 10440 2752
rect 10376 2692 10380 2748
rect 10380 2692 10436 2748
rect 10436 2692 10440 2748
rect 10376 2688 10440 2692
rect 10456 2748 10520 2752
rect 10456 2692 10460 2748
rect 10460 2692 10516 2748
rect 10516 2692 10520 2748
rect 10456 2688 10520 2692
rect 16216 2748 16280 2752
rect 16216 2692 16220 2748
rect 16220 2692 16276 2748
rect 16276 2692 16280 2748
rect 16216 2688 16280 2692
rect 16296 2748 16360 2752
rect 16296 2692 16300 2748
rect 16300 2692 16356 2748
rect 16356 2692 16360 2748
rect 16296 2688 16360 2692
rect 16376 2748 16440 2752
rect 16376 2692 16380 2748
rect 16380 2692 16436 2748
rect 16436 2692 16440 2748
rect 16376 2688 16440 2692
rect 16456 2748 16520 2752
rect 16456 2692 16460 2748
rect 16460 2692 16516 2748
rect 16516 2692 16520 2748
rect 16456 2688 16520 2692
rect 7216 2204 7280 2208
rect 7216 2148 7220 2204
rect 7220 2148 7276 2204
rect 7276 2148 7280 2204
rect 7216 2144 7280 2148
rect 7296 2204 7360 2208
rect 7296 2148 7300 2204
rect 7300 2148 7356 2204
rect 7356 2148 7360 2204
rect 7296 2144 7360 2148
rect 7376 2204 7440 2208
rect 7376 2148 7380 2204
rect 7380 2148 7436 2204
rect 7436 2148 7440 2204
rect 7376 2144 7440 2148
rect 7456 2204 7520 2208
rect 7456 2148 7460 2204
rect 7460 2148 7516 2204
rect 7516 2148 7520 2204
rect 7456 2144 7520 2148
rect 13216 2204 13280 2208
rect 13216 2148 13220 2204
rect 13220 2148 13276 2204
rect 13276 2148 13280 2204
rect 13216 2144 13280 2148
rect 13296 2204 13360 2208
rect 13296 2148 13300 2204
rect 13300 2148 13356 2204
rect 13356 2148 13360 2204
rect 13296 2144 13360 2148
rect 13376 2204 13440 2208
rect 13376 2148 13380 2204
rect 13380 2148 13436 2204
rect 13436 2148 13440 2204
rect 13376 2144 13440 2148
rect 13456 2204 13520 2208
rect 13456 2148 13460 2204
rect 13460 2148 13516 2204
rect 13516 2148 13520 2204
rect 13456 2144 13520 2148
<< metal4 >>
rect 4208 17984 4528 18000
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 7208 17440 7528 18000
rect 7208 17376 7216 17440
rect 7280 17376 7296 17440
rect 7360 17376 7376 17440
rect 7440 17376 7456 17440
rect 7520 17376 7528 17440
rect 7208 16352 7528 17376
rect 7208 16288 7216 16352
rect 7280 16288 7296 16352
rect 7360 16288 7376 16352
rect 7440 16288 7456 16352
rect 7520 16288 7528 16352
rect 7208 15264 7528 16288
rect 7208 15200 7216 15264
rect 7280 15200 7296 15264
rect 7360 15200 7376 15264
rect 7440 15200 7456 15264
rect 7520 15200 7528 15264
rect 7208 14176 7528 15200
rect 7208 14112 7216 14176
rect 7280 14112 7296 14176
rect 7360 14112 7376 14176
rect 7440 14112 7456 14176
rect 7520 14112 7528 14176
rect 7208 13088 7528 14112
rect 7208 13024 7216 13088
rect 7280 13024 7296 13088
rect 7360 13024 7376 13088
rect 7440 13024 7456 13088
rect 7520 13024 7528 13088
rect 7208 12000 7528 13024
rect 7208 11936 7216 12000
rect 7280 11936 7296 12000
rect 7360 11936 7376 12000
rect 7440 11936 7456 12000
rect 7520 11936 7528 12000
rect 7208 10912 7528 11936
rect 7208 10848 7216 10912
rect 7280 10848 7296 10912
rect 7360 10848 7376 10912
rect 7440 10848 7456 10912
rect 7520 10848 7528 10912
rect 7208 9824 7528 10848
rect 7208 9760 7216 9824
rect 7280 9760 7296 9824
rect 7360 9760 7376 9824
rect 7440 9760 7456 9824
rect 7520 9760 7528 9824
rect 7208 8736 7528 9760
rect 7208 8672 7216 8736
rect 7280 8672 7296 8736
rect 7360 8672 7376 8736
rect 7440 8672 7456 8736
rect 7520 8672 7528 8736
rect 7208 7648 7528 8672
rect 7208 7584 7216 7648
rect 7280 7584 7296 7648
rect 7360 7584 7376 7648
rect 7440 7584 7456 7648
rect 7520 7584 7528 7648
rect 7208 6560 7528 7584
rect 7208 6496 7216 6560
rect 7280 6496 7296 6560
rect 7360 6496 7376 6560
rect 7440 6496 7456 6560
rect 7520 6496 7528 6560
rect 7208 5472 7528 6496
rect 7208 5408 7216 5472
rect 7280 5408 7296 5472
rect 7360 5408 7376 5472
rect 7440 5408 7456 5472
rect 7520 5408 7528 5472
rect 7208 4384 7528 5408
rect 7208 4320 7216 4384
rect 7280 4320 7296 4384
rect 7360 4320 7376 4384
rect 7440 4320 7456 4384
rect 7520 4320 7528 4384
rect 7208 3296 7528 4320
rect 7208 3232 7216 3296
rect 7280 3232 7296 3296
rect 7360 3232 7376 3296
rect 7440 3232 7456 3296
rect 7520 3232 7528 3296
rect 7208 2208 7528 3232
rect 7208 2144 7216 2208
rect 7280 2144 7296 2208
rect 7360 2144 7376 2208
rect 7440 2144 7456 2208
rect 7520 2144 7528 2208
rect 7208 2128 7528 2144
rect 10208 17984 10528 18000
rect 10208 17920 10216 17984
rect 10280 17920 10296 17984
rect 10360 17920 10376 17984
rect 10440 17920 10456 17984
rect 10520 17920 10528 17984
rect 10208 16896 10528 17920
rect 10208 16832 10216 16896
rect 10280 16832 10296 16896
rect 10360 16832 10376 16896
rect 10440 16832 10456 16896
rect 10520 16832 10528 16896
rect 10208 15808 10528 16832
rect 10208 15744 10216 15808
rect 10280 15744 10296 15808
rect 10360 15744 10376 15808
rect 10440 15744 10456 15808
rect 10520 15744 10528 15808
rect 10208 14720 10528 15744
rect 10208 14656 10216 14720
rect 10280 14656 10296 14720
rect 10360 14656 10376 14720
rect 10440 14656 10456 14720
rect 10520 14656 10528 14720
rect 10208 13632 10528 14656
rect 10208 13568 10216 13632
rect 10280 13568 10296 13632
rect 10360 13568 10376 13632
rect 10440 13568 10456 13632
rect 10520 13568 10528 13632
rect 10208 12544 10528 13568
rect 10208 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10528 12544
rect 10208 11456 10528 12480
rect 10208 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10528 11456
rect 10208 10368 10528 11392
rect 10208 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10528 10368
rect 10208 9280 10528 10304
rect 10208 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10528 9280
rect 10208 8192 10528 9216
rect 10208 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10528 8192
rect 10208 7104 10528 8128
rect 10208 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10528 7104
rect 10208 6016 10528 7040
rect 10208 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10528 6016
rect 10208 4928 10528 5952
rect 10208 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10528 4928
rect 10208 3840 10528 4864
rect 10208 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10528 3840
rect 10208 2752 10528 3776
rect 10208 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10528 2752
rect 10208 2128 10528 2688
rect 13208 17440 13528 18000
rect 13208 17376 13216 17440
rect 13280 17376 13296 17440
rect 13360 17376 13376 17440
rect 13440 17376 13456 17440
rect 13520 17376 13528 17440
rect 13208 16352 13528 17376
rect 13208 16288 13216 16352
rect 13280 16288 13296 16352
rect 13360 16288 13376 16352
rect 13440 16288 13456 16352
rect 13520 16288 13528 16352
rect 13208 15264 13528 16288
rect 13208 15200 13216 15264
rect 13280 15200 13296 15264
rect 13360 15200 13376 15264
rect 13440 15200 13456 15264
rect 13520 15200 13528 15264
rect 13208 14176 13528 15200
rect 13208 14112 13216 14176
rect 13280 14112 13296 14176
rect 13360 14112 13376 14176
rect 13440 14112 13456 14176
rect 13520 14112 13528 14176
rect 13208 13088 13528 14112
rect 13208 13024 13216 13088
rect 13280 13024 13296 13088
rect 13360 13024 13376 13088
rect 13440 13024 13456 13088
rect 13520 13024 13528 13088
rect 13208 12000 13528 13024
rect 13208 11936 13216 12000
rect 13280 11936 13296 12000
rect 13360 11936 13376 12000
rect 13440 11936 13456 12000
rect 13520 11936 13528 12000
rect 13208 10912 13528 11936
rect 13208 10848 13216 10912
rect 13280 10848 13296 10912
rect 13360 10848 13376 10912
rect 13440 10848 13456 10912
rect 13520 10848 13528 10912
rect 13208 9824 13528 10848
rect 13208 9760 13216 9824
rect 13280 9760 13296 9824
rect 13360 9760 13376 9824
rect 13440 9760 13456 9824
rect 13520 9760 13528 9824
rect 13208 8736 13528 9760
rect 13208 8672 13216 8736
rect 13280 8672 13296 8736
rect 13360 8672 13376 8736
rect 13440 8672 13456 8736
rect 13520 8672 13528 8736
rect 13208 7648 13528 8672
rect 13208 7584 13216 7648
rect 13280 7584 13296 7648
rect 13360 7584 13376 7648
rect 13440 7584 13456 7648
rect 13520 7584 13528 7648
rect 13208 6560 13528 7584
rect 13208 6496 13216 6560
rect 13280 6496 13296 6560
rect 13360 6496 13376 6560
rect 13440 6496 13456 6560
rect 13520 6496 13528 6560
rect 13208 5472 13528 6496
rect 13208 5408 13216 5472
rect 13280 5408 13296 5472
rect 13360 5408 13376 5472
rect 13440 5408 13456 5472
rect 13520 5408 13528 5472
rect 13208 4384 13528 5408
rect 13208 4320 13216 4384
rect 13280 4320 13296 4384
rect 13360 4320 13376 4384
rect 13440 4320 13456 4384
rect 13520 4320 13528 4384
rect 13208 3296 13528 4320
rect 13208 3232 13216 3296
rect 13280 3232 13296 3296
rect 13360 3232 13376 3296
rect 13440 3232 13456 3296
rect 13520 3232 13528 3296
rect 13208 2208 13528 3232
rect 13208 2144 13216 2208
rect 13280 2144 13296 2208
rect 13360 2144 13376 2208
rect 13440 2144 13456 2208
rect 13520 2144 13528 2208
rect 13208 2128 13528 2144
rect 16208 17984 16528 18000
rect 16208 17920 16216 17984
rect 16280 17920 16296 17984
rect 16360 17920 16376 17984
rect 16440 17920 16456 17984
rect 16520 17920 16528 17984
rect 16208 16896 16528 17920
rect 16208 16832 16216 16896
rect 16280 16832 16296 16896
rect 16360 16832 16376 16896
rect 16440 16832 16456 16896
rect 16520 16832 16528 16896
rect 16208 15808 16528 16832
rect 16208 15744 16216 15808
rect 16280 15744 16296 15808
rect 16360 15744 16376 15808
rect 16440 15744 16456 15808
rect 16520 15744 16528 15808
rect 16208 14720 16528 15744
rect 16208 14656 16216 14720
rect 16280 14656 16296 14720
rect 16360 14656 16376 14720
rect 16440 14656 16456 14720
rect 16520 14656 16528 14720
rect 16208 13632 16528 14656
rect 16208 13568 16216 13632
rect 16280 13568 16296 13632
rect 16360 13568 16376 13632
rect 16440 13568 16456 13632
rect 16520 13568 16528 13632
rect 16208 12544 16528 13568
rect 16208 12480 16216 12544
rect 16280 12480 16296 12544
rect 16360 12480 16376 12544
rect 16440 12480 16456 12544
rect 16520 12480 16528 12544
rect 16208 11456 16528 12480
rect 16208 11392 16216 11456
rect 16280 11392 16296 11456
rect 16360 11392 16376 11456
rect 16440 11392 16456 11456
rect 16520 11392 16528 11456
rect 16208 10368 16528 11392
rect 16208 10304 16216 10368
rect 16280 10304 16296 10368
rect 16360 10304 16376 10368
rect 16440 10304 16456 10368
rect 16520 10304 16528 10368
rect 16208 9280 16528 10304
rect 16208 9216 16216 9280
rect 16280 9216 16296 9280
rect 16360 9216 16376 9280
rect 16440 9216 16456 9280
rect 16520 9216 16528 9280
rect 16208 8192 16528 9216
rect 16208 8128 16216 8192
rect 16280 8128 16296 8192
rect 16360 8128 16376 8192
rect 16440 8128 16456 8192
rect 16520 8128 16528 8192
rect 16208 7104 16528 8128
rect 16208 7040 16216 7104
rect 16280 7040 16296 7104
rect 16360 7040 16376 7104
rect 16440 7040 16456 7104
rect 16520 7040 16528 7104
rect 16208 6016 16528 7040
rect 16208 5952 16216 6016
rect 16280 5952 16296 6016
rect 16360 5952 16376 6016
rect 16440 5952 16456 6016
rect 16520 5952 16528 6016
rect 16208 4928 16528 5952
rect 16208 4864 16216 4928
rect 16280 4864 16296 4928
rect 16360 4864 16376 4928
rect 16440 4864 16456 4928
rect 16520 4864 16528 4928
rect 16208 3840 16528 4864
rect 16208 3776 16216 3840
rect 16280 3776 16296 3840
rect 16360 3776 16376 3840
rect 16440 3776 16456 3840
rect 16520 3776 16528 3840
rect 16208 2752 16528 3776
rect 16208 2688 16216 2752
rect 16280 2688 16296 2752
rect 16360 2688 16376 2752
rect 16440 2688 16456 2752
rect 16520 2688 16528 2752
rect 16208 2128 16528 2688
use sky130_fd_sc_hd__inv_2  _123_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 8004 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1692646696
transform -1 0 6348 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1692646696
transform -1 0 4324 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 13984 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 7360 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1692646696
transform 1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _130_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 8832 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 1692646696
transform 1 0 10028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _132_
timestamp 1692646696
transform -1 0 13156 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _133_
timestamp 1692646696
transform -1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _134_
timestamp 1692646696
transform -1 0 10212 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 1692646696
transform -1 0 5060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1692646696
transform -1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _137_
timestamp 1692646696
transform 1 0 1932 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 2576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1692646696
transform -1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _140_
timestamp 1692646696
transform 1 0 4048 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1692646696
transform 1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1692646696
transform -1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _143_
timestamp 1692646696
transform 1 0 6532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _144_
timestamp 1692646696
transform 1 0 10764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp 1692646696
transform 1 0 11684 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 11500 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 11316 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _149_
timestamp 1692646696
transform 1 0 6992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _150_
timestamp 1692646696
transform -1 0 6992 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1692646696
transform 1 0 6624 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _152_
timestamp 1692646696
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _153_
timestamp 1692646696
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1692646696
transform 1 0 6900 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _155_
timestamp 1692646696
transform 1 0 2300 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1692646696
transform 1 0 2668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _157_
timestamp 1692646696
transform 1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _158_
timestamp 1692646696
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1692646696
transform 1 0 9476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _160_
timestamp 1692646696
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _161_
timestamp 1692646696
transform 1 0 13340 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1692646696
transform 1 0 13524 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _163_
timestamp 1692646696
transform 1 0 11316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _164_
timestamp 1692646696
transform 1 0 10212 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1692646696
transform -1 0 11040 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _166_
timestamp 1692646696
transform -1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1692646696
transform -1 0 14352 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _168_
timestamp 1692646696
transform 1 0 12880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _169_
timestamp 1692646696
transform 1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _170_
timestamp 1692646696
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1692646696
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _172_
timestamp 1692646696
transform -1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _173_
timestamp 1692646696
transform -1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 10856 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _175_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 13524 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 13892 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _177_
timestamp 1692646696
transform -1 0 13248 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _178_
timestamp 1692646696
transform 1 0 13340 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _179_
timestamp 1692646696
transform -1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _180_
timestamp 1692646696
transform 1 0 13524 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _181_
timestamp 1692646696
transform 1 0 14904 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _182_
timestamp 1692646696
transform 1 0 15088 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _183_
timestamp 1692646696
transform -1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _184_
timestamp 1692646696
transform 1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 15732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 16008 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _187_
timestamp 1692646696
transform -1 0 15456 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1692646696
transform 1 0 14628 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 15180 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _190_
timestamp 1692646696
transform -1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _191_
timestamp 1692646696
transform -1 0 6808 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _192_
timestamp 1692646696
transform -1 0 6256 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1692646696
transform 1 0 5520 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _194_
timestamp 1692646696
transform -1 0 5888 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _195_
timestamp 1692646696
transform 1 0 4324 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _196_
timestamp 1692646696
transform 1 0 5520 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _197_
timestamp 1692646696
transform -1 0 5520 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _198_
timestamp 1692646696
transform -1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 5612 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _200_
timestamp 1692646696
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _201_
timestamp 1692646696
transform 1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 1692646696
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _203_
timestamp 1692646696
transform 1 0 7636 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _204_
timestamp 1692646696
transform -1 0 8556 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1692646696
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _206_
timestamp 1692646696
transform 1 0 7912 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _207_
timestamp 1692646696
transform -1 0 8740 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 7452 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _209_
timestamp 1692646696
transform -1 0 7820 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1692646696
transform -1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _211_
timestamp 1692646696
transform -1 0 8188 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 10120 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _214_
timestamp 1692646696
transform -1 0 9752 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 1692646696
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _216_
timestamp 1692646696
transform 1 0 10488 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _217_
timestamp 1692646696
transform -1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1692646696
transform -1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _220_
timestamp 1692646696
transform -1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _221_
timestamp 1692646696
transform -1 0 14812 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 14352 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 9660 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1692646696
transform -1 0 14536 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _225_
timestamp 1692646696
transform -1 0 13984 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _226_
timestamp 1692646696
transform -1 0 12696 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _227_
timestamp 1692646696
transform -1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 14720 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _229_
timestamp 1692646696
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _230_
timestamp 1692646696
transform 1 0 14076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _231_
timestamp 1692646696
transform -1 0 13432 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _232_
timestamp 1692646696
transform -1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _233_
timestamp 1692646696
transform 1 0 13432 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _234_
timestamp 1692646696
transform 1 0 12236 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 1692646696
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _236_
timestamp 1692646696
transform -1 0 11500 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 1692646696
transform 1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _238_
timestamp 1692646696
transform 1 0 11868 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _239_
timestamp 1692646696
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _240_
timestamp 1692646696
transform 1 0 11132 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _241_
timestamp 1692646696
transform 1 0 11500 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1692646696
transform 1 0 11132 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1692646696
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _244_
timestamp 1692646696
transform -1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _245_
timestamp 1692646696
transform 1 0 11960 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _246_
timestamp 1692646696
transform 1 0 11960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _247_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 12512 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _248_
timestamp 1692646696
transform 1 0 13064 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _249_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp 1692646696
transform -1 0 11408 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1692646696
transform -1 0 11684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _252_
timestamp 1692646696
transform 1 0 4048 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _253_
timestamp 1692646696
transform 1 0 4692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 1692646696
transform 1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 1692646696
transform 1 0 7084 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1692646696
transform 1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 1692646696
transform 1 0 7636 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _258_
timestamp 1692646696
transform 1 0 2760 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1692646696
transform 1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1692646696
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1692646696
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1692646696
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1692646696
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1692646696
transform 1 0 14168 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1692646696
transform -1 0 15548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1692646696
transform -1 0 14352 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _267_
timestamp 1692646696
transform -1 0 2300 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 13892 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _269_
timestamp 1692646696
transform 1 0 14904 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _270_
timestamp 1692646696
transform 1 0 14720 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _271_
timestamp 1692646696
transform -1 0 15916 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 1692646696
transform 1 0 11500 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _273_
timestamp 1692646696
transform 1 0 9568 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _274_
timestamp 1692646696
transform 1 0 9292 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _275_
timestamp 1692646696
transform 1 0 10120 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _276_
timestamp 1692646696
transform 1 0 11960 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 11500 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 1692646696
transform 1 0 4140 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _279_
timestamp 1692646696
transform 1 0 5704 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _280_
timestamp 1692646696
transform 1 0 7820 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _281_
timestamp 1692646696
transform 1 0 3496 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _282_
timestamp 1692646696
transform 1 0 4692 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _283_
timestamp 1692646696
transform 1 0 5336 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _284_
timestamp 1692646696
transform 1 0 4876 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _285_
timestamp 1692646696
transform 1 0 6624 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _286_
timestamp 1692646696
transform -1 0 9568 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _287_
timestamp 1692646696
transform 1 0 7084 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _288_
timestamp 1692646696
transform 1 0 7360 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _289_
timestamp 1692646696
transform 1 0 9476 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _290_
timestamp 1692646696
transform 1 0 6348 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _291_
timestamp 1692646696
transform 1 0 4784 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _292_
timestamp 1692646696
transform 1 0 4692 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _293_
timestamp 1692646696
transform 1 0 11684 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _294_
timestamp 1692646696
transform 1 0 9844 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _295_
timestamp 1692646696
transform 1 0 9476 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _296_
timestamp 1692646696
transform 1 0 7636 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _297_
timestamp 1692646696
transform 1 0 7360 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _298_
timestamp 1692646696
transform 1 0 6256 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _299_
timestamp 1692646696
transform 1 0 8096 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _300_
timestamp 1692646696
transform 1 0 6900 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _301_
timestamp 1692646696
transform 1 0 7820 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _302_
timestamp 1692646696
transform 1 0 6624 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _303_
timestamp 1692646696
transform 1 0 4692 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _304_
timestamp 1692646696
transform 1 0 3404 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _305_
timestamp 1692646696
transform 1 0 1748 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _306_
timestamp 1692646696
transform 1 0 2760 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _307_
timestamp 1692646696
transform 1 0 2392 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _308_
timestamp 1692646696
transform 1 0 3772 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 14076 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _309__16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 13248 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _310_
timestamp 1692646696
transform -1 0 16560 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _311_
timestamp 1692646696
transform -1 0 16560 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _312_
timestamp 1692646696
transform 1 0 5520 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _313_
timestamp 1692646696
transform 1 0 6900 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _314_
timestamp 1692646696
transform 1 0 8924 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 1692646696
transform -1 0 11408 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 1692646696
transform 1 0 11500 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _317_
timestamp 1692646696
transform 1 0 11684 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _318_
timestamp 1692646696
transform 1 0 13248 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _319_
timestamp 1692646696
transform -1 0 16192 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1692646696
transform 1 0 9108 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1692646696
transform 1 0 10488 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1692646696
transform 1 0 11500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _323_
timestamp 1692646696
transform -1 0 13892 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _324_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 7084 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _325_
timestamp 1692646696
transform 1 0 11500 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _326_
timestamp 1692646696
transform 1 0 12420 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _327_
timestamp 1692646696
transform 1 0 12972 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _328_
timestamp 1692646696
transform 1 0 14996 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _329_
timestamp 1692646696
transform -1 0 16008 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _330_
timestamp 1692646696
transform 1 0 13984 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _331_
timestamp 1692646696
transform 1 0 15272 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _332_
timestamp 1692646696
transform 1 0 14352 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1692646696
transform -1 0 16836 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _334_
timestamp 1692646696
transform 1 0 11960 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _335_
timestamp 1692646696
transform 1 0 13156 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _336_
timestamp 1692646696
transform 1 0 1564 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _337_
timestamp 1692646696
transform 1 0 2760 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _338_
timestamp 1692646696
transform 1 0 1840 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 1692646696
transform 1 0 2852 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _341_
timestamp 1692646696
transform -1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _342_
timestamp 1692646696
transform -1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _343_
timestamp 1692646696
transform -1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _344_
timestamp 1692646696
transform -1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _345_
timestamp 1692646696
transform -1 0 9200 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _346_
timestamp 1692646696
transform -1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _347_
timestamp 1692646696
transform -1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _348_
timestamp 1692646696
transform -1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _349_
timestamp 1692646696
transform -1 0 8096 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _350_
timestamp 1692646696
transform -1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _351_
timestamp 1692646696
transform -1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _352_
timestamp 1692646696
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _353_
timestamp 1692646696
transform -1 0 5060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _354_
timestamp 1692646696
transform -1 0 1932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _355_
timestamp 1692646696
transform -1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _356_
timestamp 1692646696
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _357_
timestamp 1692646696
transform -1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _358_
timestamp 1692646696
transform -1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _359_
timestamp 1692646696
transform -1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _360_
timestamp 1692646696
transform -1 0 4048 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1692646696
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__CLK
timestamp 1692646696
transform 1 0 13432 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__CLK
timestamp 1692646696
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__CLK
timestamp 1692646696
transform 1 0 14720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__CLK
timestamp 1692646696
transform 1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__CLK
timestamp 1692646696
transform -1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__CLK
timestamp 1692646696
transform -1 0 9568 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__CLK
timestamp 1692646696
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__CLK
timestamp 1692646696
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__CLK
timestamp 1692646696
transform 1 0 11776 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__CLK
timestamp 1692646696
transform 1 0 11316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__CLK
timestamp 1692646696
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__CLK
timestamp 1692646696
transform 1 0 5520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__CLK
timestamp 1692646696
transform 1 0 7636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__CLK
timestamp 1692646696
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__CLK
timestamp 1692646696
transform 1 0 4508 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__CLK
timestamp 1692646696
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__CLK
timestamp 1692646696
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__CLK
timestamp 1692646696
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__CLK
timestamp 1692646696
transform -1 0 7912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__CLK
timestamp 1692646696
transform 1 0 6900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__288__CLK
timestamp 1692646696
transform 1 0 7176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__289__CLK
timestamp 1692646696
transform 1 0 9292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__312__CLK
timestamp 1692646696
transform -1 0 4784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__324__CLK
timestamp 1692646696
transform 1 0 6900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__CLK
timestamp 1692646696
transform -1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__326__CLK
timestamp 1692646696
transform 1 0 12236 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__327__CLK
timestamp 1692646696
transform 1 0 12512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__328__CLK
timestamp 1692646696
transform 1 0 14812 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__329__CLK
timestamp 1692646696
transform 1 0 14260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__330__CLK
timestamp 1692646696
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__331__CLK
timestamp 1692646696
transform 1 0 15088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_4  fanout11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 13156 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1692646696
transform -1 0 14352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1692646696
transform -1 0 9844 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1692646696
transform 1 0 12788 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 1692646696
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1692646696
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1692646696
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_42
timestamp 1692646696
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1692646696
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1692646696
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1692646696
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1692646696
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_92
timestamp 1692646696
transform 1 0 9568 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1692646696
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1692646696
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1692646696
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_117
timestamp 1692646696
transform 1 0 11868 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_129
timestamp 1692646696
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1692646696
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1692646696
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1692646696
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_169
timestamp 1692646696
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 1692646696
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_16
timestamp 1692646696
transform 1 0 2576 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_28
timestamp 1692646696
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_40
timestamp 1692646696
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_52
timestamp 1692646696
transform 1 0 5888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_133
timestamp 1692646696
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_140
timestamp 1692646696
transform 1 0 13984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1692646696
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1692646696
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1692646696
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1692646696
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1692646696
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1692646696
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1692646696
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_37
timestamp 1692646696
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_60
timestamp 1692646696
transform 1 0 6624 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_68
timestamp 1692646696
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1692646696
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_97
timestamp 1692646696
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_105
timestamp 1692646696
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_116
timestamp 1692646696
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_120
timestamp 1692646696
transform 1 0 12144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1692646696
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_148
timestamp 1692646696
transform 1 0 14720 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_160
timestamp 1692646696
transform 1 0 15824 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_168
timestamp 1692646696
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1692646696
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_15
timestamp 1692646696
transform 1 0 2484 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_34
timestamp 1692646696
transform 1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_46
timestamp 1692646696
transform 1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_60
timestamp 1692646696
transform 1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_65
timestamp 1692646696
transform 1 0 7084 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_83
timestamp 1692646696
transform 1 0 8740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_95
timestamp 1692646696
transform 1 0 9844 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_103
timestamp 1692646696
transform 1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1692646696
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1692646696
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_128
timestamp 1692646696
transform 1 0 12880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_169
timestamp 1692646696
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1692646696
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1692646696
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1692646696
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_29
timestamp 1692646696
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_35
timestamp 1692646696
transform 1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_62
timestamp 1692646696
transform 1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1692646696
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 1692646696
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_136
timestamp 1692646696
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_146
timestamp 1692646696
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_150
timestamp 1692646696
transform 1 0 14904 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_162
timestamp 1692646696
transform 1 0 16008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_170
timestamp 1692646696
transform 1 0 16744 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1692646696
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_18
timestamp 1692646696
transform 1 0 2760 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_42
timestamp 1692646696
transform 1 0 4968 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 1692646696
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_57
timestamp 1692646696
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_63
timestamp 1692646696
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1692646696
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_105
timestamp 1692646696
transform 1 0 10764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_120
timestamp 1692646696
transform 1 0 12144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_126
timestamp 1692646696
transform 1 0 12696 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_134
timestamp 1692646696
transform 1 0 13432 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_152
timestamp 1692646696
transform 1 0 15088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_164
timestamp 1692646696
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1692646696
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1692646696
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_10
timestamp 1692646696
transform 1 0 2024 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_16
timestamp 1692646696
transform 1 0 2576 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_29
timestamp 1692646696
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_42
timestamp 1692646696
transform 1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_46
timestamp 1692646696
transform 1 0 5336 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_58
timestamp 1692646696
transform 1 0 6440 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_70
timestamp 1692646696
transform 1 0 7544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_73
timestamp 1692646696
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1692646696
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 1692646696
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_118
timestamp 1692646696
transform 1 0 11960 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_129
timestamp 1692646696
transform 1 0 12972 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_137
timestamp 1692646696
transform 1 0 13708 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_170
timestamp 1692646696
transform 1 0 16744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1692646696
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_13
timestamp 1692646696
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_32
timestamp 1692646696
transform 1 0 4048 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_36
timestamp 1692646696
transform 1 0 4416 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1692646696
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1692646696
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_65
timestamp 1692646696
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_84
timestamp 1692646696
transform 1 0 8832 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_98
timestamp 1692646696
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_102
timestamp 1692646696
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 1692646696
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1692646696
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 1692646696
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_121
timestamp 1692646696
transform 1 0 12236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_133
timestamp 1692646696
transform 1 0 13340 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_159
timestamp 1692646696
transform 1 0 15732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1692646696
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_169
timestamp 1692646696
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1692646696
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1692646696
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1692646696
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1692646696
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 1692646696
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_47
timestamp 1692646696
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1692646696
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1692646696
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_129
timestamp 1692646696
transform 1 0 12972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1692646696
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1692646696
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1692646696
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_165
timestamp 1692646696
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1692646696
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_15
timestamp 1692646696
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_19
timestamp 1692646696
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_28
timestamp 1692646696
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1692646696
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1692646696
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1692646696
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_81
timestamp 1692646696
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_97
timestamp 1692646696
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 1692646696
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1692646696
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_144
timestamp 1692646696
transform 1 0 14352 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_169
timestamp 1692646696
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_3
timestamp 1692646696
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_10
timestamp 1692646696
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_16
timestamp 1692646696
transform 1 0 2576 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1692646696
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1692646696
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1692646696
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_53
timestamp 1692646696
transform 1 0 5980 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_59
timestamp 1692646696
transform 1 0 6532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1692646696
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_85
timestamp 1692646696
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_107
timestamp 1692646696
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_111
timestamp 1692646696
transform 1 0 11316 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_115
timestamp 1692646696
transform 1 0 11684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_127
timestamp 1692646696
transform 1 0 12788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_162
timestamp 1692646696
transform 1 0 16008 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_170
timestamp 1692646696
transform 1 0 16744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1692646696
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_10
timestamp 1692646696
transform 1 0 2024 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_22
timestamp 1692646696
transform 1 0 3128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_45
timestamp 1692646696
transform 1 0 5244 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1692646696
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_66
timestamp 1692646696
transform 1 0 7176 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_72
timestamp 1692646696
transform 1 0 7728 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1692646696
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_105
timestamp 1692646696
transform 1 0 10764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_138
timestamp 1692646696
transform 1 0 13800 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 1692646696
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1692646696
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_9
timestamp 1692646696
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_13
timestamp 1692646696
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1692646696
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_29
timestamp 1692646696
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_35
timestamp 1692646696
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_67
timestamp 1692646696
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_74
timestamp 1692646696
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1692646696
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_85
timestamp 1692646696
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_89
timestamp 1692646696
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_93
timestamp 1692646696
transform 1 0 9660 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_105
timestamp 1692646696
transform 1 0 10764 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_113
timestamp 1692646696
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_125
timestamp 1692646696
transform 1 0 12604 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_131
timestamp 1692646696
transform 1 0 13156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_164
timestamp 1692646696
transform 1 0 16192 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_170
timestamp 1692646696
transform 1 0 16744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1692646696
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_7
timestamp 1692646696
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_11
timestamp 1692646696
transform 1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_17
timestamp 1692646696
transform 1 0 2668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_38
timestamp 1692646696
transform 1 0 4600 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_43
timestamp 1692646696
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1692646696
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1692646696
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_69
timestamp 1692646696
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1692646696
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1692646696
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_118
timestamp 1692646696
transform 1 0 11960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_126
timestamp 1692646696
transform 1 0 12696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_157
timestamp 1692646696
transform 1 0 15548 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1692646696
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_169
timestamp 1692646696
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_3
timestamp 1692646696
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_29
timestamp 1692646696
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_40
timestamp 1692646696
transform 1 0 4784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_51
timestamp 1692646696
transform 1 0 5796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1692646696
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1692646696
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1692646696
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_97
timestamp 1692646696
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_116
timestamp 1692646696
transform 1 0 11776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1692646696
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_147
timestamp 1692646696
transform 1 0 14628 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_9
timestamp 1692646696
transform 1 0 1932 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_17
timestamp 1692646696
transform 1 0 2668 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_26
timestamp 1692646696
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_38
timestamp 1692646696
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_62
timestamp 1692646696
transform 1 0 6808 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_70
timestamp 1692646696
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_75
timestamp 1692646696
transform 1 0 8004 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_96
timestamp 1692646696
transform 1 0 9936 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1692646696
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1692646696
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_125
timestamp 1692646696
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_144
timestamp 1692646696
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_148
timestamp 1692646696
transform 1 0 14720 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_157
timestamp 1692646696
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1692646696
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1692646696
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 1692646696
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_11
timestamp 1692646696
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_17
timestamp 1692646696
transform 1 0 2668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_25
timestamp 1692646696
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_29
timestamp 1692646696
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_40
timestamp 1692646696
transform 1 0 4784 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_48
timestamp 1692646696
transform 1 0 5520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_59
timestamp 1692646696
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1692646696
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1692646696
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_93
timestamp 1692646696
transform 1 0 9660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1692646696
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_141
timestamp 1692646696
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_149
timestamp 1692646696
transform 1 0 14812 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_157
timestamp 1692646696
transform 1 0 15548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_169
timestamp 1692646696
transform 1 0 16652 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1692646696
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_15
timestamp 1692646696
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_47
timestamp 1692646696
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1692646696
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_57
timestamp 1692646696
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_63
timestamp 1692646696
transform 1 0 6900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_67
timestamp 1692646696
transform 1 0 7268 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_75
timestamp 1692646696
transform 1 0 8004 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_87
timestamp 1692646696
transform 1 0 9108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_95
timestamp 1692646696
transform 1 0 9844 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_103
timestamp 1692646696
transform 1 0 10580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1692646696
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_113
timestamp 1692646696
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_121
timestamp 1692646696
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_146
timestamp 1692646696
transform 1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1692646696
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1692646696
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1692646696
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1692646696
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_37
timestamp 1692646696
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_55
timestamp 1692646696
transform 1 0 6164 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_59
timestamp 1692646696
transform 1 0 6532 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_63
timestamp 1692646696
transform 1 0 6900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_75
timestamp 1692646696
transform 1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1692646696
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1692646696
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_97
timestamp 1692646696
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_101
timestamp 1692646696
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_125
timestamp 1692646696
transform 1 0 12604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1692646696
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_165
timestamp 1692646696
transform 1 0 16284 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_3
timestamp 1692646696
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_9
timestamp 1692646696
transform 1 0 1932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_15
timestamp 1692646696
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_23
timestamp 1692646696
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_35
timestamp 1692646696
transform 1 0 4324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_39
timestamp 1692646696
transform 1 0 4692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_43
timestamp 1692646696
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 1692646696
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_57
timestamp 1692646696
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_64
timestamp 1692646696
transform 1 0 6992 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_108
timestamp 1692646696
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_133
timestamp 1692646696
transform 1 0 13340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_141
timestamp 1692646696
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_145
timestamp 1692646696
transform 1 0 14444 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_151
timestamp 1692646696
transform 1 0 14996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_157
timestamp 1692646696
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1692646696
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_3
timestamp 1692646696
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_9
timestamp 1692646696
transform 1 0 1932 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_21
timestamp 1692646696
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1692646696
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1692646696
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_53
timestamp 1692646696
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_76
timestamp 1692646696
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1692646696
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_107
timestamp 1692646696
transform 1 0 10948 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1692646696
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_141
timestamp 1692646696
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_150
timestamp 1692646696
transform 1 0 14904 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_159
timestamp 1692646696
transform 1 0 15732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_3
timestamp 1692646696
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_7
timestamp 1692646696
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_11
timestamp 1692646696
transform 1 0 2116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_23
timestamp 1692646696
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_37
timestamp 1692646696
transform 1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_43
timestamp 1692646696
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1692646696
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1692646696
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_69
timestamp 1692646696
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_75
timestamp 1692646696
transform 1 0 8004 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_87
timestamp 1692646696
transform 1 0 9108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_95
timestamp 1692646696
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_100
timestamp 1692646696
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1692646696
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_125
timestamp 1692646696
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_132
timestamp 1692646696
transform 1 0 13248 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_162
timestamp 1692646696
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 1692646696
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1692646696
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1692646696
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1692646696
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1692646696
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_39
timestamp 1692646696
transform 1 0 4692 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_51
timestamp 1692646696
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1692646696
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_105
timestamp 1692646696
transform 1 0 10764 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_113
timestamp 1692646696
transform 1 0 11500 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp 1692646696
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_149
timestamp 1692646696
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_3
timestamp 1692646696
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_16
timestamp 1692646696
transform 1 0 2576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_38
timestamp 1692646696
transform 1 0 4600 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_43
timestamp 1692646696
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_49
timestamp 1692646696
transform 1 0 5612 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_53
timestamp 1692646696
transform 1 0 5980 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1692646696
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_83
timestamp 1692646696
transform 1 0 8740 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_139
timestamp 1692646696
transform 1 0 13892 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_151
timestamp 1692646696
transform 1 0 14996 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_160
timestamp 1692646696
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_169
timestamp 1692646696
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 1692646696
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1692646696
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1692646696
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_37
timestamp 1692646696
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_68
timestamp 1692646696
transform 1 0 7360 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_76
timestamp 1692646696
transform 1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_94
timestamp 1692646696
transform 1 0 9752 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_98
timestamp 1692646696
transform 1 0 10120 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_110
timestamp 1692646696
transform 1 0 11224 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_113
timestamp 1692646696
transform 1 0 11500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_125
timestamp 1692646696
transform 1 0 12604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1692646696
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1692646696
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_164
timestamp 1692646696
transform 1 0 16192 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_170
timestamp 1692646696
transform 1 0 16744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_13
timestamp 1692646696
transform 1 0 2300 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_20
timestamp 1692646696
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_32
timestamp 1692646696
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_44
timestamp 1692646696
transform 1 0 5152 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1692646696
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_60
timestamp 1692646696
transform 1 0 6624 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_72
timestamp 1692646696
transform 1 0 7728 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_84
timestamp 1692646696
transform 1 0 8832 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_96
timestamp 1692646696
transform 1 0 9936 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_108
timestamp 1692646696
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1692646696
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_121
timestamp 1692646696
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_131
timestamp 1692646696
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_152
timestamp 1692646696
transform 1 0 15088 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 1692646696
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 1692646696
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 1692646696
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_11
timestamp 1692646696
transform 1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_22
timestamp 1692646696
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1692646696
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1692646696
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1692646696
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1692646696
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1692646696
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1692646696
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_109
timestamp 1692646696
transform 1 0 11132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_114
timestamp 1692646696
transform 1 0 11592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1692646696
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1692646696
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_145
timestamp 1692646696
transform 1 0 14444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_157
timestamp 1692646696
transform 1 0 15548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_169
timestamp 1692646696
transform 1 0 16652 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 1692646696
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_12
timestamp 1692646696
transform 1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_34
timestamp 1692646696
transform 1 0 4232 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_46
timestamp 1692646696
transform 1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1692646696
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_69
timestamp 1692646696
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_76
timestamp 1692646696
transform 1 0 8096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_84
timestamp 1692646696
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_88
timestamp 1692646696
transform 1 0 9200 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_100
timestamp 1692646696
transform 1 0 10304 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_105
timestamp 1692646696
transform 1 0 10764 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_139
timestamp 1692646696
transform 1 0 13892 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_151
timestamp 1692646696
transform 1 0 14996 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_163
timestamp 1692646696
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1692646696
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_169
timestamp 1692646696
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_6
timestamp 1692646696
transform 1 0 1656 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_14
timestamp 1692646696
transform 1 0 2392 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_20
timestamp 1692646696
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1692646696
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1692646696
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_53
timestamp 1692646696
transform 1 0 5980 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_57
timestamp 1692646696
transform 1 0 6348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_69
timestamp 1692646696
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1692646696
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1692646696
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1692646696
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_109
timestamp 1692646696
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_113
timestamp 1692646696
transform 1 0 11500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_125
timestamp 1692646696
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1692646696
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1692646696
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_153
timestamp 1692646696
transform 1 0 15180 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_167
timestamp 1692646696
transform 1 0 16468 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_169
timestamp 1692646696
transform 1 0 16652 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1692646696
transform -1 0 14076 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1692646696
transform 1 0 13892 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1692646696
transform -1 0 16560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1692646696
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1692646696
transform -1 0 16192 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1692646696
transform -1 0 16468 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1692646696
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1692646696
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1692646696
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1692646696
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  MS_CLK_RST_17
timestamp 1692646696
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output9
timestamp 1692646696
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1692646696
transform -1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_29
timestamp 1692646696
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1692646696
transform -1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_30
timestamp 1692646696
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1692646696
transform -1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_31
timestamp 1692646696
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1692646696
transform -1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_32
timestamp 1692646696
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1692646696
transform -1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_33
timestamp 1692646696
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1692646696
transform -1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_34
timestamp 1692646696
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1692646696
transform -1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_35
timestamp 1692646696
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1692646696
transform -1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_36
timestamp 1692646696
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1692646696
transform -1 0 17112 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_37
timestamp 1692646696
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1692646696
transform -1 0 17112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_38
timestamp 1692646696
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1692646696
transform -1 0 17112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_39
timestamp 1692646696
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1692646696
transform -1 0 17112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_40
timestamp 1692646696
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1692646696
transform -1 0 17112 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_41
timestamp 1692646696
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1692646696
transform -1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_42
timestamp 1692646696
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1692646696
transform -1 0 17112 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_43
timestamp 1692646696
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1692646696
transform -1 0 17112 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_44
timestamp 1692646696
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1692646696
transform -1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_45
timestamp 1692646696
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1692646696
transform -1 0 17112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_46
timestamp 1692646696
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1692646696
transform -1 0 17112 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_47
timestamp 1692646696
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1692646696
transform -1 0 17112 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_48
timestamp 1692646696
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1692646696
transform -1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_49
timestamp 1692646696
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1692646696
transform -1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_50
timestamp 1692646696
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1692646696
transform -1 0 17112 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_51
timestamp 1692646696
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1692646696
transform -1 0 17112 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_52
timestamp 1692646696
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1692646696
transform -1 0 17112 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_53
timestamp 1692646696
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1692646696
transform -1 0 17112 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_54
timestamp 1692646696
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1692646696
transform -1 0 17112 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_55
timestamp 1692646696
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1692646696
transform -1 0 17112 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_56
timestamp 1692646696
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1692646696
transform -1 0 17112 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_57
timestamp 1692646696
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1692646696
transform -1 0 17112 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  PoR.ROSC_CLKBUF_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 2668 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  PoR.ROSC_CLKBUF_1
timestamp 1692646696
transform 1 0 3220 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYBUF_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 2944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_0.clkdlybuf
timestamp 1692646696
transform -1 0 6256 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_0.clkinv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 10764 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_1.clkdlybuf
timestamp 1692646696
transform -1 0 5980 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_1.clkinv
timestamp 1692646696
transform 1 0 5612 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_2.clkdlybuf
timestamp 1692646696
transform -1 0 5520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_2.clkinv
timestamp 1692646696
transform -1 0 5612 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_3.clkdlybuf
timestamp 1692646696
transform -1 0 4692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_3.clkinv
timestamp 1692646696
transform -1 0 5060 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_4.clkdlybuf
timestamp 1692646696
transform -1 0 4140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_4.clkinv
timestamp 1692646696
transform 1 0 4140 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_5.clkdlybuf
timestamp 1692646696
transform -1 0 3496 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_5.clkinv
timestamp 1692646696
transform -1 0 3680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  PoR.ROSC_DLYINV_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform -1 0 3772 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1692646696
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1692646696
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1692646696
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1692646696
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 1692646696
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 1692646696
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 1692646696
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_65
timestamp 1692646696
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_66
timestamp 1692646696
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 1692646696
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_68
timestamp 1692646696
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_69
timestamp 1692646696
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 1692646696
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_71
timestamp 1692646696
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_72
timestamp 1692646696
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 1692646696
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_74
timestamp 1692646696
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp 1692646696
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 1692646696
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp 1692646696
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp 1692646696
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 1692646696
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp 1692646696
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp 1692646696
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1692646696
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp 1692646696
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp 1692646696
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 1692646696
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_86
timestamp 1692646696
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp 1692646696
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 1692646696
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp 1692646696
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_90
timestamp 1692646696
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 1692646696
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp 1692646696
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp 1692646696
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 1692646696
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_95
timestamp 1692646696
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp 1692646696
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 1692646696
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_98
timestamp 1692646696
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_99
timestamp 1692646696
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 1692646696
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_101
timestamp 1692646696
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_102
timestamp 1692646696
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 1692646696
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_104
timestamp 1692646696
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_105
timestamp 1692646696
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 1692646696
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_107
timestamp 1692646696
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_108
timestamp 1692646696
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 1692646696
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_110
timestamp 1692646696
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_111
timestamp 1692646696
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 1692646696
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_113
timestamp 1692646696
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_114
timestamp 1692646696
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 1692646696
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_116
timestamp 1692646696
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_117
timestamp 1692646696
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 1692646696
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_119
timestamp 1692646696
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_120
timestamp 1692646696
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 1692646696
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_122
timestamp 1692646696
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_123
timestamp 1692646696
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 1692646696
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_125
timestamp 1692646696
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_126
timestamp 1692646696
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 1692646696
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_128
timestamp 1692646696
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_129
timestamp 1692646696
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 1692646696
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_131
timestamp 1692646696
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_132
timestamp 1692646696
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 1692646696
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_134
timestamp 1692646696
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_135
timestamp 1692646696
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 1692646696
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_137
timestamp 1692646696
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_138
timestamp 1692646696
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 1692646696
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_140
timestamp 1692646696
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_141
timestamp 1692646696
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 1692646696
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 1692646696
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 1692646696
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_145
timestamp 1692646696
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_146
timestamp 1692646696
transform 1 0 6256 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_147
timestamp 1692646696
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_148
timestamp 1692646696
transform 1 0 11408 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 1692646696
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 1692646696
transform 1 0 16560 0 1 17408
box -38 -48 130 592
<< labels >>
flabel metal3 s 17506 12248 18306 12368 0 FreeSans 480 0 0 0 clk
port 0 nsew signal tristate
flabel metal2 s 5814 19650 5870 20450 0 FreeSans 224 90 0 0 clk_div[0]
port 1 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 clk_div[1]
port 2 nsew signal input
flabel metal2 s 10966 19650 11022 20450 0 FreeSans 224 90 0 0 por_fb_in
port 3 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 por_fb_out
port 4 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 por_n
port 5 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 rst_n
port 6 nsew signal tristate
flabel metal3 s 17506 1368 18306 1488 0 FreeSans 480 0 0 0 sel_mux0
port 7 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 sel_mux1
port 8 nsew signal input
flabel metal3 s 17506 17688 18306 17808 0 FreeSans 480 0 0 0 sel_mux2
port 9 nsew signal input
flabel metal2 s 16118 19650 16174 20450 0 FreeSans 224 90 0 0 sel_rosc[0]
port 10 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 sel_rosc[1]
port 11 nsew signal input
flabel metal4 s 4208 2128 4528 18000 0 FreeSans 1920 90 0 0 vccd1
port 12 nsew power bidirectional
flabel metal4 s 10208 2128 10528 18000 0 FreeSans 1920 90 0 0 vccd1
port 12 nsew power bidirectional
flabel metal4 s 16208 2128 16528 18000 0 FreeSans 1920 90 0 0 vccd1
port 12 nsew power bidirectional
flabel metal4 s 7208 2128 7528 18000 0 FreeSans 1920 90 0 0 vssd1
port 13 nsew ground bidirectional
flabel metal4 s 13208 2128 13528 18000 0 FreeSans 1920 90 0 0 vssd1
port 13 nsew ground bidirectional
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 xclk0
port 14 nsew signal input
flabel metal2 s 662 19650 718 20450 0 FreeSans 224 90 0 0 xclk1
port 15 nsew signal input
flabel metal3 s 17506 6808 18306 6928 0 FreeSans 480 0 0 0 xrst_n
port 16 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 18306 20450
<< end >>
