magic
tech sky130A
magscale 1 2
timestamp 1694343306
<< viali >>
rect 7113 21573 7147 21607
rect 14197 21573 14231 21607
rect 3801 21505 3835 21539
rect 6929 21505 6963 21539
rect 7389 21505 7423 21539
rect 7573 21505 7607 21539
rect 10333 21505 10367 21539
rect 18981 21505 19015 21539
rect 20269 21505 20303 21539
rect 4077 21437 4111 21471
rect 10057 21437 10091 21471
rect 10885 21437 10919 21471
rect 7297 21301 7331 21335
rect 7481 21301 7515 21335
rect 14289 21301 14323 21335
rect 18797 21301 18831 21335
rect 20361 21301 20395 21335
rect 7665 21097 7699 21131
rect 5917 20961 5951 20995
rect 6285 20961 6319 20995
rect 8217 20961 8251 20995
rect 4721 20893 4755 20927
rect 6009 20893 6043 20927
rect 8033 20893 8067 20927
rect 9597 20893 9631 20927
rect 10333 20893 10367 20927
rect 10600 20893 10634 20927
rect 13921 20893 13955 20927
rect 16497 20893 16531 20927
rect 6530 20825 6564 20859
rect 7849 20825 7883 20859
rect 8585 20825 8619 20859
rect 13654 20825 13688 20859
rect 16764 20825 16798 20859
rect 4537 20757 4571 20791
rect 6193 20757 6227 20791
rect 9413 20757 9447 20791
rect 10149 20757 10183 20791
rect 11713 20757 11747 20791
rect 12541 20757 12575 20791
rect 17877 20757 17911 20791
rect 8493 20553 8527 20587
rect 18490 20485 18524 20519
rect 4537 20417 4571 20451
rect 13470 20417 13504 20451
rect 13737 20417 13771 20451
rect 15873 20417 15907 20451
rect 17886 20417 17920 20451
rect 6745 20349 6779 20383
rect 7021 20349 7055 20383
rect 10057 20349 10091 20383
rect 10333 20349 10367 20383
rect 16129 20349 16163 20383
rect 18153 20349 18187 20383
rect 18245 20349 18279 20383
rect 3893 20213 3927 20247
rect 6653 20213 6687 20247
rect 8585 20213 8619 20247
rect 12357 20213 12391 20247
rect 14749 20213 14783 20247
rect 16773 20213 16807 20247
rect 19625 20213 19659 20247
rect 6009 20009 6043 20043
rect 8401 20009 8435 20043
rect 10241 20009 10275 20043
rect 13553 20009 13587 20043
rect 14105 20009 14139 20043
rect 6377 19941 6411 19975
rect 6469 19873 6503 19907
rect 9781 19873 9815 19907
rect 3893 19805 3927 19839
rect 6101 19805 6135 19839
rect 7113 19805 7147 19839
rect 7205 19805 7239 19839
rect 7389 19805 7423 19839
rect 8493 19805 8527 19839
rect 8953 19805 8987 19839
rect 9597 19805 9631 19839
rect 9873 19805 9907 19839
rect 12173 19805 12207 19839
rect 12440 19805 12474 19839
rect 14105 19805 14139 19839
rect 14197 19805 14231 19839
rect 15393 19805 15427 19839
rect 15649 19805 15683 19839
rect 17233 19805 17267 19839
rect 19073 19805 19107 19839
rect 6377 19737 6411 19771
rect 16957 19737 16991 19771
rect 18828 19737 18862 19771
rect 3893 19669 3927 19703
rect 6193 19669 6227 19703
rect 7297 19669 7331 19703
rect 14473 19669 14507 19703
rect 16773 19669 16807 19703
rect 17141 19669 17175 19703
rect 17325 19669 17359 19703
rect 17509 19669 17543 19703
rect 17693 19669 17727 19703
rect 4629 19465 4663 19499
rect 6469 19465 6503 19499
rect 10149 19465 10183 19499
rect 11805 19465 11839 19499
rect 13369 19465 13403 19499
rect 16129 19465 16163 19499
rect 4261 19397 4295 19431
rect 7582 19397 7616 19431
rect 9321 19397 9355 19431
rect 13537 19397 13571 19431
rect 13737 19397 13771 19431
rect 16681 19397 16715 19431
rect 2513 19329 2547 19363
rect 3157 19329 3191 19363
rect 3249 19329 3283 19363
rect 3985 19329 4019 19363
rect 4721 19329 4755 19363
rect 4988 19329 5022 19363
rect 9045 19329 9079 19363
rect 9229 19329 9263 19363
rect 10057 19329 10091 19363
rect 10333 19329 10367 19363
rect 10517 19329 10551 19363
rect 13277 19329 13311 19363
rect 16497 19329 16531 19363
rect 18788 19329 18822 19363
rect 3893 19261 3927 19295
rect 7849 19261 7883 19295
rect 9873 19261 9907 19295
rect 11161 19261 11195 19295
rect 16405 19261 16439 19295
rect 18521 19261 18555 19295
rect 6101 19193 6135 19227
rect 9045 19125 9079 19159
rect 10333 19125 10367 19159
rect 13553 19125 13587 19159
rect 16497 19125 16531 19159
rect 17969 19125 18003 19159
rect 19901 19125 19935 19159
rect 5089 18921 5123 18955
rect 6653 18921 6687 18955
rect 6837 18921 6871 18955
rect 8769 18921 8803 18955
rect 9229 18921 9263 18955
rect 11253 18921 11287 18955
rect 16681 18921 16715 18955
rect 16865 18921 16899 18955
rect 17141 18921 17175 18955
rect 18981 18921 19015 18955
rect 2789 18853 2823 18887
rect 9413 18853 9447 18887
rect 20269 18853 20303 18887
rect 5733 18785 5767 18819
rect 5825 18785 5859 18819
rect 6101 18785 6135 18819
rect 7021 18785 7055 18819
rect 11621 18785 11655 18819
rect 17601 18785 17635 18819
rect 2697 18717 2731 18751
rect 2789 18717 2823 18751
rect 6193 18717 6227 18751
rect 9505 18717 9539 18751
rect 11888 18717 11922 18751
rect 15301 18717 15335 18751
rect 15568 18717 15602 18751
rect 17049 18717 17083 18751
rect 17141 18717 17175 18751
rect 17325 18717 17359 18751
rect 17857 18717 17891 18751
rect 20085 18717 20119 18751
rect 6469 18649 6503 18683
rect 6669 18649 6703 18683
rect 7297 18649 7331 18683
rect 9045 18649 9079 18683
rect 9781 18649 9815 18683
rect 19993 18649 20027 18683
rect 2053 18581 2087 18615
rect 9255 18581 9289 18615
rect 13001 18581 13035 18615
rect 19717 18581 19751 18615
rect 19901 18581 19935 18615
rect 6929 18377 6963 18411
rect 8861 18377 8895 18411
rect 9229 18377 9263 18411
rect 9321 18377 9355 18411
rect 9781 18377 9815 18411
rect 15393 18377 15427 18411
rect 16681 18377 16715 18411
rect 17693 18377 17727 18411
rect 9597 18309 9631 18343
rect 13654 18309 13688 18343
rect 14280 18309 14314 18343
rect 17233 18309 17267 18343
rect 17449 18309 17483 18343
rect 17861 18309 17895 18343
rect 18061 18309 18095 18343
rect 18880 18309 18914 18343
rect 2145 18241 2179 18275
rect 8769 18241 8803 18275
rect 8953 18241 8987 18275
rect 9045 18241 9079 18275
rect 9413 18241 9447 18275
rect 9689 18241 9723 18275
rect 9873 18241 9907 18275
rect 13921 18241 13955 18275
rect 14013 18241 14047 18275
rect 16865 18241 16899 18275
rect 17049 18241 17083 18275
rect 18613 18241 18647 18275
rect 2145 18037 2179 18071
rect 10241 18037 10275 18071
rect 12541 18037 12575 18071
rect 16865 18037 16899 18071
rect 17417 18037 17451 18071
rect 17601 18037 17635 18071
rect 17877 18037 17911 18071
rect 19993 18037 20027 18071
rect 14749 17833 14783 17867
rect 19257 17833 19291 17867
rect 19625 17833 19659 17867
rect 17785 17765 17819 17799
rect 5273 17697 5307 17731
rect 16129 17697 16163 17731
rect 17877 17697 17911 17731
rect 19625 17697 19659 17731
rect 3249 17629 3283 17663
rect 3801 17629 3835 17663
rect 4445 17629 4479 17663
rect 4537 17629 4571 17663
rect 4721 17629 4755 17663
rect 4905 17629 4939 17663
rect 5089 17629 5123 17663
rect 5365 17629 5399 17663
rect 5549 17629 5583 17663
rect 9965 17629 9999 17663
rect 13001 17629 13035 17663
rect 15862 17629 15896 17663
rect 17601 17629 17635 17663
rect 19441 17629 19475 17663
rect 19717 17629 19751 17663
rect 2982 17561 3016 17595
rect 10232 17561 10266 17595
rect 12734 17561 12768 17595
rect 13093 17561 13127 17595
rect 13369 17561 13403 17595
rect 13461 17561 13495 17595
rect 17969 17561 18003 17595
rect 1869 17493 1903 17527
rect 3617 17493 3651 17527
rect 4629 17493 4663 17527
rect 5457 17493 5491 17527
rect 5641 17493 5675 17527
rect 11345 17493 11379 17527
rect 11621 17493 11655 17527
rect 13277 17493 13311 17527
rect 13645 17493 13679 17527
rect 17693 17493 17727 17527
rect 1685 17289 1719 17323
rect 2697 17289 2731 17323
rect 17049 17289 17083 17323
rect 4016 17221 4050 17255
rect 13277 17221 13311 17255
rect 13493 17221 13527 17255
rect 1777 17153 1811 17187
rect 6837 17153 6871 17187
rect 9321 17153 9355 17187
rect 10241 17153 10275 17187
rect 12633 17153 12667 17187
rect 12909 17153 12943 17187
rect 13737 17153 13771 17187
rect 18173 17153 18207 17187
rect 19248 17153 19282 17187
rect 1869 17085 1903 17119
rect 2053 17085 2087 17119
rect 4261 17085 4295 17119
rect 4353 17085 4387 17119
rect 4629 17085 4663 17119
rect 7113 17085 7147 17119
rect 9413 17085 9447 17119
rect 10885 17085 10919 17119
rect 12725 17085 12759 17119
rect 13829 17085 13863 17119
rect 18429 17085 18463 17119
rect 18981 17085 19015 17119
rect 13093 17017 13127 17051
rect 2881 16949 2915 16983
rect 6101 16949 6135 16983
rect 8585 16949 8619 16983
rect 9597 16949 9631 16983
rect 12909 16949 12943 16983
rect 13461 16949 13495 16983
rect 13645 16949 13679 16983
rect 13829 16949 13863 16983
rect 14105 16949 14139 16983
rect 20361 16949 20395 16983
rect 3985 16745 4019 16779
rect 6180 16745 6214 16779
rect 7665 16745 7699 16779
rect 11069 16745 11103 16779
rect 18613 16745 18647 16779
rect 19073 16745 19107 16779
rect 14933 16677 14967 16711
rect 19809 16677 19843 16711
rect 1685 16609 1719 16643
rect 5825 16609 5859 16643
rect 9321 16609 9355 16643
rect 9597 16609 9631 16643
rect 15117 16609 15151 16643
rect 15209 16609 15243 16643
rect 15485 16609 15519 16643
rect 15577 16609 15611 16643
rect 15761 16609 15795 16643
rect 16037 16609 16071 16643
rect 17877 16609 17911 16643
rect 18061 16609 18095 16643
rect 3341 16541 3375 16575
rect 5917 16541 5951 16575
rect 8493 16541 8527 16575
rect 8585 16541 8619 16575
rect 8769 16541 8803 16575
rect 9137 16541 9171 16575
rect 11161 16541 11195 16575
rect 11428 16541 11462 16575
rect 14933 16541 14967 16575
rect 15301 16541 15335 16575
rect 15393 16541 15427 16575
rect 15853 16541 15887 16575
rect 17785 16541 17819 16575
rect 18153 16541 18187 16575
rect 18797 16541 18831 16575
rect 18889 16541 18923 16575
rect 19533 16541 19567 16575
rect 1501 16473 1535 16507
rect 3074 16473 3108 16507
rect 3801 16473 3835 16507
rect 5558 16473 5592 16507
rect 17601 16473 17635 16507
rect 18245 16473 18279 16507
rect 19073 16473 19107 16507
rect 19441 16473 19475 16507
rect 1961 16405 1995 16439
rect 4001 16405 4035 16439
rect 4169 16405 4203 16439
rect 4445 16405 4479 16439
rect 8217 16405 8251 16439
rect 8953 16405 8987 16439
rect 12541 16405 12575 16439
rect 19257 16405 19291 16439
rect 19625 16405 19659 16439
rect 2697 16201 2731 16235
rect 3249 16201 3283 16235
rect 4261 16201 4295 16235
rect 9597 16201 9631 16235
rect 9689 16201 9723 16235
rect 10149 16201 10183 16235
rect 14933 16201 14967 16235
rect 16773 16201 16807 16235
rect 19993 16201 20027 16235
rect 3433 16133 3467 16167
rect 3617 16133 3651 16167
rect 4997 16133 5031 16167
rect 8125 16133 8159 16167
rect 9873 16133 9907 16167
rect 18880 16133 18914 16167
rect 1593 16065 1627 16099
rect 3341 16065 3375 16099
rect 4905 16065 4939 16099
rect 5089 16065 5123 16099
rect 10057 16065 10091 16099
rect 10149 16065 10183 16099
rect 10333 16065 10367 16099
rect 13165 16065 13199 16099
rect 14473 16065 14507 16099
rect 14749 16065 14783 16099
rect 15281 16065 15315 16099
rect 17886 16065 17920 16099
rect 18153 16065 18187 16099
rect 18613 16065 18647 16099
rect 1685 15997 1719 16031
rect 1961 15997 1995 16031
rect 2053 15997 2087 16031
rect 7849 15997 7883 16031
rect 12909 15997 12943 16031
rect 14657 15997 14691 16031
rect 15025 15997 15059 16031
rect 3617 15929 3651 15963
rect 16405 15929 16439 15963
rect 7757 15861 7791 15895
rect 14289 15861 14323 15895
rect 14749 15861 14783 15895
rect 13461 15657 13495 15691
rect 13921 15657 13955 15691
rect 15669 15657 15703 15691
rect 6837 15589 6871 15623
rect 12817 15589 12851 15623
rect 13369 15589 13403 15623
rect 16221 15589 16255 15623
rect 6929 15521 6963 15555
rect 11253 15521 11287 15555
rect 2053 15453 2087 15487
rect 4169 15453 4203 15487
rect 7205 15453 7239 15487
rect 13001 15453 13035 15487
rect 13093 15453 13127 15487
rect 13645 15453 13679 15487
rect 13737 15453 13771 15487
rect 14105 15453 14139 15487
rect 14372 15453 14406 15487
rect 15853 15453 15887 15487
rect 17325 15453 17359 15487
rect 17509 15453 17543 15487
rect 17693 15453 17727 15487
rect 17785 15453 17819 15487
rect 18061 15453 18095 15487
rect 6469 15385 6503 15419
rect 11520 15385 11554 15419
rect 13461 15385 13495 15419
rect 15945 15385 15979 15419
rect 17141 15385 17175 15419
rect 1961 15317 1995 15351
rect 4261 15317 4295 15351
rect 7021 15317 7055 15351
rect 12633 15317 12667 15351
rect 13185 15317 13219 15351
rect 15485 15317 15519 15351
rect 16037 15317 16071 15351
rect 17417 15317 17451 15351
rect 9873 15113 9907 15147
rect 13185 15113 13219 15147
rect 15577 15113 15611 15147
rect 19901 15113 19935 15147
rect 3801 15045 3835 15079
rect 3893 15045 3927 15079
rect 6653 15045 6687 15079
rect 9965 15045 9999 15079
rect 14464 15045 14498 15079
rect 18788 15045 18822 15079
rect 1409 14977 1443 15011
rect 3341 14977 3375 15011
rect 3617 14977 3651 15011
rect 3985 14977 4019 15011
rect 10057 14977 10091 15011
rect 10609 14977 10643 15011
rect 10793 14977 10827 15011
rect 11805 14977 11839 15011
rect 12072 14977 12106 15011
rect 18521 14977 18555 15011
rect 1685 14909 1719 14943
rect 4261 14909 4295 14943
rect 5733 14909 5767 14943
rect 6009 14909 6043 14943
rect 6377 14909 6411 14943
rect 10517 14909 10551 14943
rect 10701 14909 10735 14943
rect 14197 14909 14231 14943
rect 10241 14841 10275 14875
rect 3157 14773 3191 14807
rect 3525 14773 3559 14807
rect 4169 14773 4203 14807
rect 8125 14773 8159 14807
rect 8953 14773 8987 14807
rect 9689 14773 9723 14807
rect 10333 14773 10367 14807
rect 1593 14569 1627 14603
rect 3617 14569 3651 14603
rect 10793 14569 10827 14603
rect 11437 14569 11471 14603
rect 17141 14569 17175 14603
rect 2145 14433 2179 14467
rect 7297 14433 7331 14467
rect 9045 14433 9079 14467
rect 12817 14433 12851 14467
rect 15301 14433 15335 14467
rect 16957 14433 16991 14467
rect 17601 14433 17635 14467
rect 1593 14365 1627 14399
rect 1777 14365 1811 14399
rect 1869 14365 1903 14399
rect 7021 14365 7055 14399
rect 12550 14365 12584 14399
rect 17134 14365 17168 14399
rect 5181 14297 5215 14331
rect 6929 14297 6963 14331
rect 9321 14297 9355 14331
rect 15568 14297 15602 14331
rect 16865 14297 16899 14331
rect 17846 14297 17880 14331
rect 8769 14229 8803 14263
rect 16681 14229 16715 14263
rect 17325 14229 17359 14263
rect 18981 14229 19015 14263
rect 3249 14025 3283 14059
rect 5549 14025 5583 14059
rect 5825 14025 5859 14059
rect 7665 14025 7699 14059
rect 9965 14025 9999 14059
rect 11805 14025 11839 14059
rect 18153 14025 18187 14059
rect 4077 13957 4111 13991
rect 8585 13957 8619 13991
rect 8677 13957 8711 13991
rect 9413 13957 9447 13991
rect 14565 13957 14599 13991
rect 16313 13957 16347 13991
rect 16681 13957 16715 13991
rect 18880 13957 18914 13991
rect 3709 13889 3743 13923
rect 3801 13889 3835 13923
rect 5733 13889 5767 13923
rect 6009 13889 6043 13923
rect 6193 13889 6227 13923
rect 6377 13889 6411 13923
rect 8441 13889 8475 13923
rect 8861 13889 8895 13923
rect 10149 13889 10183 13923
rect 13277 13889 13311 13923
rect 9873 13821 9907 13855
rect 18613 13821 18647 13855
rect 3341 13753 3375 13787
rect 9781 13753 9815 13787
rect 6009 13685 6043 13719
rect 8309 13685 8343 13719
rect 10517 13685 10551 13719
rect 19993 13685 20027 13719
rect 4800 13481 4834 13515
rect 8125 13481 8159 13515
rect 18061 13481 18095 13515
rect 15669 13413 15703 13447
rect 16497 13413 16531 13447
rect 4537 13345 4571 13379
rect 6285 13345 6319 13379
rect 6653 13345 6687 13379
rect 9781 13345 9815 13379
rect 10241 13345 10275 13379
rect 10333 13345 10367 13379
rect 13001 13345 13035 13379
rect 14289 13345 14323 13379
rect 3341 13277 3375 13311
rect 3525 13277 3559 13311
rect 4261 13277 4295 13311
rect 6377 13277 6411 13311
rect 9137 13277 9171 13311
rect 9873 13277 9907 13311
rect 13369 13277 13403 13311
rect 15945 13277 15979 13311
rect 16681 13277 16715 13311
rect 9321 13209 9355 13243
rect 10609 13209 10643 13243
rect 12173 13209 12207 13243
rect 13921 13209 13955 13243
rect 14545 13209 14579 13243
rect 16129 13209 16163 13243
rect 16221 13209 16255 13243
rect 16926 13209 16960 13243
rect 2513 13141 2547 13175
rect 3433 13141 3467 13175
rect 4169 13141 4203 13175
rect 4353 13141 4387 13175
rect 8953 13141 8987 13175
rect 12081 13141 12115 13175
rect 13553 13141 13587 13175
rect 13645 13141 13679 13175
rect 13737 13141 13771 13175
rect 16313 13141 16347 13175
rect 7021 12937 7055 12971
rect 7941 12937 7975 12971
rect 9781 12937 9815 12971
rect 10701 12937 10735 12971
rect 11621 12937 11655 12971
rect 12265 12937 12299 12971
rect 14197 12937 14231 12971
rect 16773 12937 16807 12971
rect 18705 12937 18739 12971
rect 20361 12937 20395 12971
rect 2881 12869 2915 12903
rect 10149 12869 10183 12903
rect 15310 12869 15344 12903
rect 17886 12869 17920 12903
rect 18521 12869 18555 12903
rect 1685 12801 1719 12835
rect 2605 12801 2639 12835
rect 4445 12801 4479 12835
rect 6377 12801 6411 12835
rect 6745 12801 6779 12835
rect 6929 12801 6963 12835
rect 8033 12801 8067 12835
rect 10517 12801 10551 12835
rect 11345 12801 11379 12835
rect 11897 12801 11931 12835
rect 13378 12801 13412 12835
rect 15669 12801 15703 12835
rect 15945 12801 15979 12835
rect 18153 12801 18187 12835
rect 18613 12801 18647 12835
rect 19248 12801 19282 12835
rect 2421 12733 2455 12767
rect 4353 12733 4387 12767
rect 4721 12733 4755 12767
rect 8309 12733 8343 12767
rect 13645 12733 13679 12767
rect 15577 12733 15611 12767
rect 15853 12733 15887 12767
rect 18981 12733 19015 12767
rect 2145 12665 2179 12699
rect 9965 12665 9999 12699
rect 18889 12665 18923 12699
rect 1777 12597 1811 12631
rect 1961 12597 1995 12631
rect 6193 12597 6227 12631
rect 10149 12597 10183 12631
rect 15761 12597 15795 12631
rect 16129 12597 16163 12631
rect 18337 12597 18371 12631
rect 3617 12393 3651 12427
rect 4353 12393 4387 12427
rect 8585 12393 8619 12427
rect 9321 12393 9355 12427
rect 14197 12393 14231 12427
rect 19257 12393 19291 12427
rect 20085 12393 20119 12427
rect 18981 12325 19015 12359
rect 19717 12325 19751 12359
rect 19993 12325 20027 12359
rect 17601 12257 17635 12291
rect 19441 12257 19475 12291
rect 1777 12189 1811 12223
rect 1869 12189 1903 12223
rect 3801 12189 3835 12223
rect 4221 12189 4255 12223
rect 8769 12189 8803 12223
rect 9137 12189 9171 12223
rect 9597 12189 9631 12223
rect 13277 12189 13311 12223
rect 15577 12189 15611 12223
rect 15669 12189 15703 12223
rect 17868 12189 17902 12223
rect 19257 12189 19291 12223
rect 19533 12189 19567 12223
rect 2145 12121 2179 12155
rect 3985 12121 4019 12155
rect 4077 12121 4111 12155
rect 9505 12121 9539 12155
rect 15310 12121 15344 12155
rect 15936 12121 15970 12155
rect 19809 12121 19843 12155
rect 20177 12121 20211 12155
rect 1593 12053 1627 12087
rect 12725 12053 12759 12087
rect 17049 12053 17083 12087
rect 19901 12053 19935 12087
rect 3157 11849 3191 11883
rect 3709 11849 3743 11883
rect 12173 11849 12207 11883
rect 16221 11849 16255 11883
rect 16881 11849 16915 11883
rect 17509 11849 17543 11883
rect 20361 11849 20395 11883
rect 1685 11781 1719 11815
rect 15853 11781 15887 11815
rect 16053 11781 16087 11815
rect 16681 11781 16715 11815
rect 17969 11781 18003 11815
rect 18521 11781 18555 11815
rect 19226 11781 19260 11815
rect 1409 11713 1443 11747
rect 8677 11713 8711 11747
rect 9781 11713 9815 11747
rect 11069 11713 11103 11747
rect 13297 11713 13331 11747
rect 13553 11713 13587 11747
rect 13645 11713 13679 11747
rect 17141 11713 17175 11747
rect 18153 11713 18187 11747
rect 18981 11713 19015 11747
rect 17233 11645 17267 11679
rect 18245 11645 18279 11679
rect 18429 11645 18463 11679
rect 18613 11645 18647 11679
rect 17049 11577 17083 11611
rect 8493 11509 8527 11543
rect 9965 11509 9999 11543
rect 10977 11509 11011 11543
rect 14933 11509 14967 11543
rect 16037 11509 16071 11543
rect 16865 11509 16899 11543
rect 17141 11509 17175 11543
rect 1593 11305 1627 11339
rect 5181 11305 5215 11339
rect 7665 11305 7699 11339
rect 8585 11305 8619 11339
rect 8769 11305 8803 11339
rect 12725 11305 12759 11339
rect 17601 11305 17635 11339
rect 18153 11305 18187 11339
rect 19625 11305 19659 11339
rect 18521 11237 18555 11271
rect 19257 11237 19291 11271
rect 5273 11169 5307 11203
rect 9321 11169 9355 11203
rect 10793 11169 10827 11203
rect 11161 11169 11195 11203
rect 13369 11169 13403 11203
rect 1409 11101 1443 11135
rect 9045 11101 9079 11135
rect 10885 11101 10919 11135
rect 13645 11101 13679 11135
rect 15669 11101 15703 11135
rect 18153 11101 18187 11135
rect 18245 11101 18279 11135
rect 19441 11101 19475 11135
rect 19533 11101 19567 11135
rect 5549 11033 5583 11067
rect 8217 11033 8251 11067
rect 8401 11033 8435 11067
rect 8617 11033 8651 11067
rect 13553 11033 13587 11067
rect 14105 11033 14139 11067
rect 16313 11033 16347 11067
rect 19717 11033 19751 11067
rect 7021 10965 7055 10999
rect 8125 10965 8159 10999
rect 12633 10965 12667 10999
rect 3249 10761 3283 10795
rect 5549 10761 5583 10795
rect 7481 10761 7515 10795
rect 9551 10761 9585 10795
rect 15669 10761 15703 10795
rect 16773 10761 16807 10795
rect 19993 10761 20027 10795
rect 4537 10693 4571 10727
rect 5273 10693 5307 10727
rect 10977 10693 11011 10727
rect 20177 10693 20211 10727
rect 2237 10625 2271 10659
rect 4813 10625 4847 10659
rect 4997 10625 5031 10659
rect 5457 10625 5491 10659
rect 5825 10625 5859 10659
rect 6101 10625 6135 10659
rect 6377 10625 6411 10659
rect 7021 10625 7055 10659
rect 7113 10625 7147 10659
rect 7297 10625 7331 10659
rect 7573 10625 7607 10659
rect 9965 10625 9999 10659
rect 10425 10625 10459 10659
rect 10701 10625 10735 10659
rect 10885 10625 10919 10659
rect 11121 10625 11155 10659
rect 11621 10625 11655 10659
rect 12081 10625 12115 10659
rect 13921 10625 13955 10659
rect 17886 10625 17920 10659
rect 18153 10625 18187 10659
rect 18245 10625 18279 10659
rect 18512 10625 18546 10659
rect 20085 10625 20119 10659
rect 4905 10557 4939 10591
rect 5733 10557 5767 10591
rect 6193 10557 6227 10591
rect 7757 10557 7791 10591
rect 8125 10557 8159 10591
rect 14197 10557 14231 10591
rect 10241 10489 10275 10523
rect 11253 10489 11287 10523
rect 19809 10489 19843 10523
rect 1593 10421 1627 10455
rect 5089 10421 5123 10455
rect 7113 10421 7147 10455
rect 9689 10421 9723 10455
rect 10057 10421 10091 10455
rect 10149 10421 10183 10455
rect 11713 10421 11747 10455
rect 13369 10421 13403 10455
rect 19625 10421 19659 10455
rect 20361 10421 20395 10455
rect 3617 10217 3651 10251
rect 5549 10217 5583 10251
rect 6653 10217 6687 10251
rect 8493 10217 8527 10251
rect 8953 10217 8987 10251
rect 10701 10217 10735 10251
rect 13185 10217 13219 10251
rect 15761 10217 15795 10251
rect 18429 10217 18463 10251
rect 20269 10217 20303 10251
rect 1869 10081 1903 10115
rect 6193 10081 6227 10115
rect 6745 10081 6779 10115
rect 11437 10081 11471 10115
rect 18889 10081 18923 10115
rect 3801 10013 3835 10047
rect 9321 10013 9355 10047
rect 9781 10013 9815 10047
rect 10517 10013 10551 10047
rect 10701 10013 10735 10047
rect 11161 10013 11195 10047
rect 11345 10013 11379 10047
rect 13829 10013 13863 10047
rect 14381 10013 14415 10047
rect 16773 10013 16807 10047
rect 17040 10013 17074 10047
rect 18613 10013 18647 10047
rect 18705 10013 18739 10047
rect 19073 10013 19107 10047
rect 20361 10013 20395 10047
rect 2145 9945 2179 9979
rect 4077 9945 4111 9979
rect 7021 9945 7055 9979
rect 9137 9945 9171 9979
rect 9873 9945 9907 9979
rect 11253 9945 11287 9979
rect 11713 9945 11747 9979
rect 13277 9945 13311 9979
rect 14648 9945 14682 9979
rect 18981 9945 19015 9979
rect 5641 9877 5675 9911
rect 18153 9877 18187 9911
rect 2789 9673 2823 9707
rect 6929 9673 6963 9707
rect 7481 9673 7515 9707
rect 12449 9673 12483 9707
rect 18797 9673 18831 9707
rect 4629 9605 4663 9639
rect 4997 9605 5031 9639
rect 6561 9605 6595 9639
rect 7389 9605 7423 9639
rect 9347 9605 9381 9639
rect 9965 9605 9999 9639
rect 1777 9537 1811 9571
rect 2973 9537 3007 9571
rect 4169 9537 4203 9571
rect 4813 9537 4847 9571
rect 4905 9537 4939 9571
rect 5115 9537 5149 9571
rect 5273 9537 5307 9571
rect 5641 9537 5675 9571
rect 5917 9537 5951 9571
rect 6377 9537 6411 9571
rect 6653 9537 6687 9571
rect 6745 9537 6779 9571
rect 7021 9537 7055 9571
rect 7205 9537 7239 9571
rect 7757 9537 7791 9571
rect 7849 9537 7883 9571
rect 8033 9537 8067 9571
rect 9137 9537 9171 9571
rect 9229 9537 9263 9571
rect 9597 9537 9631 9571
rect 10517 9537 10551 9571
rect 12357 9537 12391 9571
rect 12633 9537 12667 9571
rect 14473 9537 14507 9571
rect 14740 9537 14774 9571
rect 17417 9537 17451 9571
rect 17684 9537 17718 9571
rect 19248 9537 19282 9571
rect 4261 9469 4295 9503
rect 4445 9469 4479 9503
rect 5733 9469 5767 9503
rect 7481 9469 7515 9503
rect 8953 9469 8987 9503
rect 18981 9469 19015 9503
rect 3801 9401 3835 9435
rect 7665 9401 7699 9435
rect 9597 9401 9631 9435
rect 1777 9333 1811 9367
rect 3341 9333 3375 9367
rect 3709 9333 3743 9367
rect 5917 9333 5951 9367
rect 6101 9333 6135 9367
rect 7849 9333 7883 9367
rect 8401 9333 8435 9367
rect 9505 9333 9539 9367
rect 12173 9333 12207 9367
rect 15853 9333 15887 9367
rect 20361 9333 20395 9367
rect 5549 9129 5583 9163
rect 5733 9129 5767 9163
rect 6929 9129 6963 9163
rect 9229 9129 9263 9163
rect 17785 9129 17819 9163
rect 17877 9129 17911 9163
rect 18245 9129 18279 9163
rect 18429 9129 18463 9163
rect 17601 9061 17635 9095
rect 17969 8993 18003 9027
rect 1593 8925 1627 8959
rect 4813 8925 4847 8959
rect 5089 8925 5123 8959
rect 8953 8925 8987 8959
rect 9229 8925 9263 8959
rect 9505 8925 9539 8959
rect 13369 8925 13403 8959
rect 13461 8925 13495 8959
rect 16241 8925 16275 8959
rect 16497 8925 16531 8959
rect 4905 8857 4939 8891
rect 5365 8857 5399 8891
rect 5581 8857 5615 8891
rect 8309 8857 8343 8891
rect 9781 8857 9815 8891
rect 11345 8857 11379 8891
rect 13093 8857 13127 8891
rect 17601 8857 17635 8891
rect 18061 8857 18095 8891
rect 2237 8789 2271 8823
rect 4997 8789 5031 8823
rect 8401 8789 8435 8823
rect 9045 8789 9079 8823
rect 11253 8789 11287 8823
rect 13185 8789 13219 8823
rect 13553 8789 13587 8823
rect 15117 8789 15151 8823
rect 18271 8789 18305 8823
rect 5917 8585 5951 8619
rect 8033 8585 8067 8619
rect 11270 8585 11304 8619
rect 14013 8585 14047 8619
rect 16405 8585 16439 8619
rect 19901 8585 19935 8619
rect 4261 8517 4295 8551
rect 4471 8517 4505 8551
rect 4721 8517 4755 8551
rect 5733 8517 5767 8551
rect 6745 8517 6779 8551
rect 6929 8517 6963 8551
rect 7129 8517 7163 8551
rect 8585 8517 8619 8551
rect 9137 8517 9171 8551
rect 10885 8517 10919 8551
rect 12541 8517 12575 8551
rect 14381 8517 14415 8551
rect 16037 8517 16071 8551
rect 16253 8517 16287 8551
rect 2421 8449 2455 8483
rect 4169 8449 4203 8483
rect 4353 8449 4387 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 5178 8449 5212 8483
rect 5549 8449 5583 8483
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 6837 8449 6871 8483
rect 7573 8449 7607 8483
rect 8861 8449 8895 8483
rect 10701 8449 10735 8483
rect 10977 8449 11011 8483
rect 11097 8449 11131 8483
rect 12265 8449 12299 8483
rect 14105 8449 14139 8483
rect 16681 8449 16715 8483
rect 18429 8449 18463 8483
rect 18521 8449 18555 8483
rect 18788 8449 18822 8483
rect 4629 8381 4663 8415
rect 6101 8381 6135 8415
rect 11621 8381 11655 8415
rect 12173 8381 12207 8415
rect 7297 8313 7331 8347
rect 8217 8313 8251 8347
rect 8769 8313 8803 8347
rect 10609 8313 10643 8347
rect 15853 8313 15887 8347
rect 1777 8245 1811 8279
rect 3985 8245 4019 8279
rect 6377 8245 6411 8279
rect 7113 8245 7147 8279
rect 7481 8245 7515 8279
rect 8585 8245 8619 8279
rect 16221 8245 16255 8279
rect 5549 8041 5583 8075
rect 9413 8041 9447 8075
rect 10793 8041 10827 8075
rect 13645 8041 13679 8075
rect 16681 8041 16715 8075
rect 17233 8041 17267 8075
rect 17509 8041 17543 8075
rect 19257 8041 19291 8075
rect 19993 8041 20027 8075
rect 6469 7973 6503 8007
rect 11713 7973 11747 8007
rect 17049 7973 17083 8007
rect 18981 7973 19015 8007
rect 19809 7973 19843 8007
rect 20361 7973 20395 8007
rect 6377 7905 6411 7939
rect 8769 7905 8803 7939
rect 17233 7905 17267 7939
rect 1777 7837 1811 7871
rect 3617 7837 3651 7871
rect 3801 7837 3835 7871
rect 5917 7837 5951 7871
rect 6101 7837 6135 7871
rect 6745 7837 6779 7871
rect 6929 7837 6963 7871
rect 10701 7837 10735 7871
rect 11345 7837 11379 7871
rect 11529 7837 11563 7871
rect 11897 7837 11931 7871
rect 15117 7837 15151 7871
rect 16681 7837 16715 7871
rect 16773 7837 16807 7871
rect 17141 7837 17175 7871
rect 17601 7837 17635 7871
rect 19533 7837 19567 7871
rect 20085 7837 20119 7871
rect 20177 7837 20211 7871
rect 2513 7769 2547 7803
rect 4077 7769 4111 7803
rect 5733 7769 5767 7803
rect 6009 7769 6043 7803
rect 6239 7769 6273 7803
rect 8493 7769 8527 7803
rect 12173 7769 12207 7803
rect 15384 7769 15418 7803
rect 17868 7769 17902 7803
rect 19901 7769 19935 7803
rect 6653 7701 6687 7735
rect 7021 7701 7055 7735
rect 16497 7701 16531 7735
rect 19441 7701 19475 7735
rect 19625 7701 19659 7735
rect 4629 7497 4663 7531
rect 5733 7497 5767 7531
rect 6377 7497 6411 7531
rect 8125 7497 8159 7531
rect 8677 7497 8711 7531
rect 12449 7497 12483 7531
rect 17233 7497 17267 7531
rect 19993 7497 20027 7531
rect 2697 7429 2731 7463
rect 4997 7429 5031 7463
rect 5365 7429 5399 7463
rect 9965 7429 9999 7463
rect 15884 7429 15918 7463
rect 18880 7429 18914 7463
rect 4813 7361 4847 7395
rect 4905 7361 4939 7395
rect 5181 7361 5215 7395
rect 5273 7361 5307 7395
rect 5457 7361 5491 7395
rect 5917 7361 5951 7395
rect 6193 7361 6227 7395
rect 6929 7361 6963 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 10701 7361 10735 7395
rect 10885 7361 10919 7395
rect 11621 7361 11655 7395
rect 11713 7361 11747 7395
rect 11897 7361 11931 7395
rect 12541 7361 12575 7395
rect 16129 7361 16163 7395
rect 16773 7361 16807 7395
rect 17049 7361 17083 7395
rect 18613 7361 18647 7395
rect 2421 7293 2455 7327
rect 4169 7293 4203 7327
rect 6101 7293 6135 7327
rect 7481 7293 7515 7327
rect 16865 7293 16899 7327
rect 10517 7225 10551 7259
rect 11161 7225 11195 7259
rect 11345 7225 11379 7259
rect 2329 7157 2363 7191
rect 5917 7157 5951 7191
rect 7389 7157 7423 7191
rect 11713 7157 11747 7191
rect 14749 7157 14783 7191
rect 16957 7157 16991 7191
rect 4800 6953 4834 6987
rect 6285 6953 6319 6987
rect 10701 6953 10735 6987
rect 18981 6953 19015 6987
rect 16773 6885 16807 6919
rect 11069 6817 11103 6851
rect 15209 6817 15243 6851
rect 17325 6817 17359 6851
rect 4537 6749 4571 6783
rect 6377 6749 6411 6783
rect 6561 6749 6595 6783
rect 6745 6749 6779 6783
rect 7573 6749 7607 6783
rect 8217 6749 8251 6783
rect 8953 6749 8987 6783
rect 10977 6749 11011 6783
rect 11161 6749 11195 6783
rect 15476 6749 15510 6783
rect 17141 6749 17175 6783
rect 17601 6749 17635 6783
rect 6653 6681 6687 6715
rect 7021 6681 7055 6715
rect 8033 6681 8067 6715
rect 8769 6681 8803 6715
rect 9229 6681 9263 6715
rect 17049 6681 17083 6715
rect 17868 6681 17902 6715
rect 4445 6613 4479 6647
rect 6929 6613 6963 6647
rect 16589 6613 16623 6647
rect 16957 6613 16991 6647
rect 6193 6409 6227 6443
rect 12541 6409 12575 6443
rect 18061 6409 18095 6443
rect 19625 6409 19659 6443
rect 2421 6341 2455 6375
rect 6653 6341 6687 6375
rect 12909 6341 12943 6375
rect 18490 6341 18524 6375
rect 2697 6273 2731 6307
rect 6377 6273 6411 6307
rect 9965 6273 9999 6307
rect 10057 6273 10091 6307
rect 10793 6273 10827 6307
rect 11529 6273 11563 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 11949 6273 11983 6307
rect 12357 6273 12391 6307
rect 16681 6273 16715 6307
rect 16948 6273 16982 6307
rect 18245 6273 18279 6307
rect 1593 6205 1627 6239
rect 2789 6205 2823 6239
rect 3065 6205 3099 6239
rect 8125 6205 8159 6239
rect 12633 6205 12667 6239
rect 14473 6205 14507 6239
rect 14749 6205 14783 6239
rect 10701 6137 10735 6171
rect 12081 6137 12115 6171
rect 14381 6137 14415 6171
rect 2513 6069 2547 6103
rect 4537 6069 4571 6103
rect 8677 6069 8711 6103
rect 10241 6069 10275 6103
rect 16221 6069 16255 6103
rect 3433 5865 3467 5899
rect 5549 5865 5583 5899
rect 7389 5865 7423 5899
rect 9045 5865 9079 5899
rect 13645 5865 13679 5899
rect 17325 5865 17359 5899
rect 13553 5797 13587 5831
rect 13737 5797 13771 5831
rect 14565 5797 14599 5831
rect 1685 5729 1719 5763
rect 1961 5729 1995 5763
rect 5641 5729 5675 5763
rect 9505 5729 9539 5763
rect 15945 5729 15979 5763
rect 1409 5661 1443 5695
rect 7481 5661 7515 5695
rect 8953 5661 8987 5695
rect 9229 5661 9263 5695
rect 9413 5661 9447 5695
rect 11345 5661 11379 5695
rect 13737 5661 13771 5695
rect 13921 5661 13955 5695
rect 15853 5661 15887 5695
rect 16212 5661 16246 5695
rect 5917 5593 5951 5627
rect 9781 5593 9815 5627
rect 13185 5593 13219 5627
rect 1593 5525 1627 5559
rect 7665 5525 7699 5559
rect 9321 5525 9355 5559
rect 11253 5525 11287 5559
rect 12633 5525 12667 5559
rect 2513 5321 2547 5355
rect 3157 5321 3191 5355
rect 4353 5321 4387 5355
rect 9229 5321 9263 5355
rect 12817 5321 12851 5355
rect 14289 5321 14323 5355
rect 14565 5321 14599 5355
rect 2329 5253 2363 5287
rect 10701 5253 10735 5287
rect 11529 5253 11563 5287
rect 14197 5253 14231 5287
rect 1501 5185 1535 5219
rect 3249 5185 3283 5219
rect 3341 5185 3375 5219
rect 3525 5185 3559 5219
rect 3801 5185 3835 5219
rect 3985 5185 4019 5219
rect 4077 5185 4111 5219
rect 4169 5185 4203 5219
rect 8493 5185 8527 5219
rect 8677 5185 8711 5219
rect 8769 5185 8803 5219
rect 8889 5185 8923 5219
rect 11253 5185 11287 5219
rect 14473 5185 14507 5219
rect 20453 5185 20487 5219
rect 2973 5117 3007 5151
rect 4445 5117 4479 5151
rect 4721 5117 4755 5151
rect 6469 5117 6503 5151
rect 10977 5117 11011 5151
rect 13921 5117 13955 5151
rect 2605 5049 2639 5083
rect 9045 5049 9079 5083
rect 3341 4981 3375 5015
rect 6193 4981 6227 5015
rect 6726 4981 6760 5015
rect 8217 4981 8251 5015
rect 11069 4981 11103 5015
rect 13369 4981 13403 5015
rect 20269 4981 20303 5015
rect 4629 4777 4663 4811
rect 5365 4777 5399 4811
rect 6377 4777 6411 4811
rect 12173 4777 12207 4811
rect 4077 4573 4111 4607
rect 4445 4573 4479 4607
rect 5273 4573 5307 4607
rect 6285 4573 6319 4607
rect 9045 4573 9079 4607
rect 13553 4573 13587 4607
rect 13645 4573 13679 4607
rect 13829 4573 13863 4607
rect 4261 4505 4295 4539
rect 4353 4505 4387 4539
rect 10885 4505 10919 4539
rect 10333 4437 10367 4471
rect 13461 4437 13495 4471
rect 13737 4437 13771 4471
rect 12909 4233 12943 4267
rect 8585 4165 8619 4199
rect 13369 4165 13403 4199
rect 3985 4097 4019 4131
rect 8033 4097 8067 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 8493 4097 8527 4131
rect 8682 4097 8716 4131
rect 9045 4097 9079 4131
rect 9229 4097 9263 4131
rect 9321 4097 9355 4131
rect 9418 4097 9452 4131
rect 10232 4097 10266 4131
rect 11529 4097 11563 4131
rect 11796 4097 11830 4131
rect 9965 4029 9999 4063
rect 13093 4029 13127 4063
rect 9597 3961 9631 3995
rect 4077 3893 4111 3927
rect 8033 3893 8067 3927
rect 8861 3893 8895 3927
rect 11345 3893 11379 3927
rect 14841 3893 14875 3927
rect 3985 3689 4019 3723
rect 9689 3689 9723 3723
rect 12541 3689 12575 3723
rect 13553 3621 13587 3655
rect 5733 3553 5767 3587
rect 7297 3553 7331 3587
rect 10241 3553 10275 3587
rect 13645 3553 13679 3587
rect 14381 3553 14415 3587
rect 7021 3485 7055 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 9557 3485 9591 3519
rect 9873 3485 9907 3519
rect 12357 3485 12391 3519
rect 12725 3485 12759 3519
rect 12817 3485 12851 3519
rect 13093 3485 13127 3519
rect 13921 3485 13955 3519
rect 14105 3485 14139 3519
rect 5457 3417 5491 3451
rect 9321 3417 9355 3451
rect 10508 3417 10542 3451
rect 12909 3417 12943 3451
rect 13185 3417 13219 3451
rect 8769 3349 8803 3383
rect 9965 3349 9999 3383
rect 11621 3349 11655 3383
rect 11805 3349 11839 3383
rect 13737 3349 13771 3383
rect 15853 3349 15887 3383
rect 5089 3145 5123 3179
rect 8493 3145 8527 3179
rect 11529 3145 11563 3179
rect 16129 3145 16163 3179
rect 3617 3077 3651 3111
rect 12817 3077 12851 3111
rect 10241 3009 10275 3043
rect 12265 3009 12299 3043
rect 12449 3009 12483 3043
rect 12541 3009 12575 3043
rect 3341 2941 3375 2975
rect 9965 2941 9999 2975
rect 10425 2941 10459 2975
rect 10701 2941 10735 2975
rect 12081 2941 12115 2975
rect 14381 2941 14415 2975
rect 14657 2941 14691 2975
rect 14289 2873 14323 2907
rect 12357 2805 12391 2839
rect 9413 2601 9447 2635
rect 11989 2601 12023 2635
rect 13277 2601 13311 2635
rect 5457 2533 5491 2567
rect 13645 2533 13679 2567
rect 7021 2465 7055 2499
rect 10977 2465 11011 2499
rect 11345 2465 11379 2499
rect 11621 2465 11655 2499
rect 5273 2397 5307 2431
rect 8769 2397 8803 2431
rect 10701 2397 10735 2431
rect 11161 2397 11195 2431
rect 11713 2397 11747 2431
rect 13185 2397 13219 2431
rect 13553 2397 13587 2431
rect 15761 2397 15795 2431
rect 12173 2329 12207 2363
rect 12357 2329 12391 2363
rect 12541 2329 12575 2363
rect 15577 2329 15611 2363
<< metal1 >>
rect 1104 21786 20792 21808
rect 1104 21734 7214 21786
rect 7266 21734 7278 21786
rect 7330 21734 7342 21786
rect 7394 21734 7406 21786
rect 7458 21734 7470 21786
rect 7522 21734 13214 21786
rect 13266 21734 13278 21786
rect 13330 21734 13342 21786
rect 13394 21734 13406 21786
rect 13458 21734 13470 21786
rect 13522 21734 19214 21786
rect 19266 21734 19278 21786
rect 19330 21734 19342 21786
rect 19394 21734 19406 21786
rect 19458 21734 19470 21786
rect 19522 21734 20792 21786
rect 1104 21712 20792 21734
rect 7101 21607 7159 21613
rect 7101 21573 7113 21607
rect 7147 21604 7159 21607
rect 7147 21576 7604 21604
rect 7147 21573 7159 21576
rect 7101 21567 7159 21573
rect 3234 21496 3240 21548
rect 3292 21536 3298 21548
rect 3789 21539 3847 21545
rect 3789 21536 3801 21539
rect 3292 21508 3801 21536
rect 3292 21496 3298 21508
rect 3789 21505 3801 21508
rect 3835 21505 3847 21539
rect 3789 21499 3847 21505
rect 6914 21496 6920 21548
rect 6972 21536 6978 21548
rect 7576 21545 7604 21576
rect 13814 21564 13820 21616
rect 13872 21604 13878 21616
rect 14185 21607 14243 21613
rect 14185 21604 14197 21607
rect 13872 21576 14197 21604
rect 13872 21564 13878 21576
rect 14185 21573 14197 21576
rect 14231 21573 14243 21607
rect 14185 21567 14243 21573
rect 7377 21539 7435 21545
rect 7377 21536 7389 21539
rect 6972 21508 7389 21536
rect 6972 21496 6978 21508
rect 7377 21505 7389 21508
rect 7423 21505 7435 21539
rect 7377 21499 7435 21505
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 10321 21539 10379 21545
rect 7607 21508 7696 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 4065 21471 4123 21477
rect 4065 21437 4077 21471
rect 4111 21468 4123 21471
rect 5718 21468 5724 21480
rect 4111 21440 5724 21468
rect 4111 21437 4123 21440
rect 4065 21431 4123 21437
rect 5718 21428 5724 21440
rect 5776 21428 5782 21480
rect 7668 21344 7696 21508
rect 10321 21505 10333 21539
rect 10367 21536 10379 21539
rect 11514 21536 11520 21548
rect 10367 21508 11520 21536
rect 10367 21505 10379 21508
rect 10321 21499 10379 21505
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 18690 21496 18696 21548
rect 18748 21536 18754 21548
rect 18969 21539 19027 21545
rect 18969 21536 18981 21539
rect 18748 21508 18981 21536
rect 18748 21496 18754 21508
rect 18969 21505 18981 21508
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 20254 21496 20260 21548
rect 20312 21496 20318 21548
rect 10042 21428 10048 21480
rect 10100 21428 10106 21480
rect 10870 21428 10876 21480
rect 10928 21428 10934 21480
rect 7282 21292 7288 21344
rect 7340 21292 7346 21344
rect 7469 21335 7527 21341
rect 7469 21301 7481 21335
rect 7515 21332 7527 21335
rect 7558 21332 7564 21344
rect 7515 21304 7564 21332
rect 7515 21301 7527 21304
rect 7469 21295 7527 21301
rect 7558 21292 7564 21304
rect 7616 21292 7622 21344
rect 7650 21292 7656 21344
rect 7708 21292 7714 21344
rect 14274 21292 14280 21344
rect 14332 21292 14338 21344
rect 18230 21292 18236 21344
rect 18288 21332 18294 21344
rect 18785 21335 18843 21341
rect 18785 21332 18797 21335
rect 18288 21304 18797 21332
rect 18288 21292 18294 21304
rect 18785 21301 18797 21304
rect 18831 21301 18843 21335
rect 18785 21295 18843 21301
rect 20349 21335 20407 21341
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20438 21332 20444 21344
rect 20395 21304 20444 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20438 21292 20444 21304
rect 20496 21292 20502 21344
rect 1104 21242 20792 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 10214 21242
rect 10266 21190 10278 21242
rect 10330 21190 10342 21242
rect 10394 21190 10406 21242
rect 10458 21190 10470 21242
rect 10522 21190 16214 21242
rect 16266 21190 16278 21242
rect 16330 21190 16342 21242
rect 16394 21190 16406 21242
rect 16458 21190 16470 21242
rect 16522 21190 20792 21242
rect 1104 21168 20792 21190
rect 5828 21100 7236 21128
rect 4709 20927 4767 20933
rect 4709 20893 4721 20927
rect 4755 20924 4767 20927
rect 5828 20924 5856 21100
rect 7208 21060 7236 21100
rect 7650 21088 7656 21140
rect 7708 21088 7714 21140
rect 8386 21088 8392 21140
rect 8444 21088 8450 21140
rect 10042 21088 10048 21140
rect 10100 21088 10106 21140
rect 8404 21060 8432 21088
rect 7208 21032 8432 21060
rect 5905 20995 5963 21001
rect 5905 20961 5917 20995
rect 5951 20992 5963 20995
rect 6270 20992 6276 21004
rect 5951 20964 6276 20992
rect 5951 20961 5963 20964
rect 5905 20955 5963 20961
rect 6270 20952 6276 20964
rect 6328 20952 6334 21004
rect 7282 20952 7288 21004
rect 7340 20952 7346 21004
rect 7558 20952 7564 21004
rect 7616 20992 7622 21004
rect 8205 20995 8263 21001
rect 8205 20992 8217 20995
rect 7616 20964 8217 20992
rect 7616 20952 7622 20964
rect 8205 20961 8217 20964
rect 8251 20992 8263 20995
rect 10060 20992 10088 21088
rect 8251 20964 10088 20992
rect 8251 20961 8263 20964
rect 8205 20955 8263 20961
rect 4755 20896 5856 20924
rect 5997 20927 6055 20933
rect 4755 20893 4767 20896
rect 4709 20887 4767 20893
rect 5997 20893 6009 20927
rect 6043 20924 6055 20927
rect 7300 20924 7328 20952
rect 8021 20927 8079 20933
rect 8021 20924 8033 20927
rect 6043 20896 6960 20924
rect 7300 20896 8033 20924
rect 6043 20893 6055 20896
rect 5997 20887 6055 20893
rect 6518 20859 6576 20865
rect 6518 20856 6530 20859
rect 6196 20828 6530 20856
rect 4522 20748 4528 20800
rect 4580 20748 4586 20800
rect 6196 20797 6224 20828
rect 6518 20825 6530 20828
rect 6564 20825 6576 20859
rect 6932 20856 6960 20896
rect 8021 20893 8033 20896
rect 8067 20893 8079 20927
rect 9582 20924 9588 20936
rect 8021 20887 8079 20893
rect 8496 20896 9588 20924
rect 7837 20859 7895 20865
rect 7837 20856 7849 20859
rect 6932 20828 7849 20856
rect 6518 20819 6576 20825
rect 7837 20825 7849 20828
rect 7883 20825 7895 20859
rect 7837 20819 7895 20825
rect 8496 20800 8524 20896
rect 9582 20884 9588 20896
rect 9640 20884 9646 20936
rect 10321 20927 10379 20933
rect 10321 20924 10333 20927
rect 10152 20896 10333 20924
rect 8573 20859 8631 20865
rect 8573 20825 8585 20859
rect 8619 20856 8631 20859
rect 8619 20828 9720 20856
rect 8619 20825 8631 20828
rect 8573 20819 8631 20825
rect 9692 20800 9720 20828
rect 6181 20791 6239 20797
rect 6181 20757 6193 20791
rect 6227 20757 6239 20791
rect 6181 20751 6239 20757
rect 8478 20748 8484 20800
rect 8536 20748 8542 20800
rect 9398 20748 9404 20800
rect 9456 20748 9462 20800
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 10152 20797 10180 20896
rect 10321 20893 10333 20896
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 10588 20927 10646 20933
rect 10588 20893 10600 20927
rect 10634 20924 10646 20927
rect 10870 20924 10876 20936
rect 10634 20896 10876 20924
rect 10634 20893 10646 20896
rect 10588 20887 10646 20893
rect 10870 20884 10876 20896
rect 10928 20884 10934 20936
rect 11716 20896 13768 20924
rect 11716 20797 11744 20896
rect 13642 20859 13700 20865
rect 13642 20825 13654 20859
rect 13688 20825 13700 20859
rect 13740 20856 13768 20896
rect 13814 20884 13820 20936
rect 13872 20924 13878 20936
rect 13909 20927 13967 20933
rect 13909 20924 13921 20927
rect 13872 20896 13921 20924
rect 13872 20884 13878 20896
rect 13909 20893 13921 20896
rect 13955 20893 13967 20927
rect 13909 20887 13967 20893
rect 16114 20884 16120 20936
rect 16172 20924 16178 20936
rect 16485 20927 16543 20933
rect 16485 20924 16497 20927
rect 16172 20896 16497 20924
rect 16172 20884 16178 20896
rect 16485 20893 16497 20896
rect 16531 20893 16543 20927
rect 16485 20887 16543 20893
rect 14550 20856 14556 20868
rect 13740 20828 14556 20856
rect 13642 20819 13700 20825
rect 10137 20791 10195 20797
rect 10137 20788 10149 20791
rect 9732 20760 10149 20788
rect 9732 20748 9738 20760
rect 10137 20757 10149 20760
rect 10183 20757 10195 20791
rect 10137 20751 10195 20757
rect 11701 20791 11759 20797
rect 11701 20757 11713 20791
rect 11747 20757 11759 20791
rect 11701 20751 11759 20757
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 12529 20791 12587 20797
rect 12529 20788 12541 20791
rect 12492 20760 12541 20788
rect 12492 20748 12498 20760
rect 12529 20757 12541 20760
rect 12575 20757 12587 20791
rect 13648 20788 13676 20819
rect 14550 20816 14556 20828
rect 14608 20816 14614 20868
rect 16752 20859 16810 20865
rect 16752 20825 16764 20859
rect 16798 20856 16810 20859
rect 17126 20856 17132 20868
rect 16798 20828 17132 20856
rect 16798 20825 16810 20828
rect 16752 20819 16810 20825
rect 17126 20816 17132 20828
rect 17184 20816 17190 20868
rect 14274 20788 14280 20800
rect 13648 20760 14280 20788
rect 12529 20751 12587 20757
rect 14274 20748 14280 20760
rect 14332 20748 14338 20800
rect 17034 20748 17040 20800
rect 17092 20788 17098 20800
rect 17862 20788 17868 20800
rect 17092 20760 17868 20788
rect 17092 20748 17098 20760
rect 17862 20748 17868 20760
rect 17920 20748 17926 20800
rect 1104 20698 20792 20720
rect 1104 20646 7214 20698
rect 7266 20646 7278 20698
rect 7330 20646 7342 20698
rect 7394 20646 7406 20698
rect 7458 20646 7470 20698
rect 7522 20646 13214 20698
rect 13266 20646 13278 20698
rect 13330 20646 13342 20698
rect 13394 20646 13406 20698
rect 13458 20646 13470 20698
rect 13522 20646 19214 20698
rect 19266 20646 19278 20698
rect 19330 20646 19342 20698
rect 19394 20646 19406 20698
rect 19458 20646 19470 20698
rect 19522 20646 20792 20698
rect 1104 20624 20792 20646
rect 8478 20544 8484 20596
rect 8536 20544 8542 20596
rect 17862 20544 17868 20596
rect 17920 20544 17926 20596
rect 8294 20516 8300 20528
rect 8234 20488 8300 20516
rect 8294 20476 8300 20488
rect 8352 20516 8358 20528
rect 8352 20488 8878 20516
rect 8352 20476 8358 20488
rect 11514 20476 11520 20528
rect 11572 20516 11578 20528
rect 13814 20516 13820 20528
rect 11572 20488 13820 20516
rect 11572 20476 11578 20488
rect 4522 20408 4528 20460
rect 4580 20408 4586 20460
rect 13446 20408 13452 20460
rect 13504 20457 13510 20460
rect 13740 20457 13768 20488
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 17880 20516 17908 20544
rect 18478 20519 18536 20525
rect 18478 20516 18490 20519
rect 17880 20488 18490 20516
rect 18478 20485 18490 20488
rect 18524 20485 18536 20519
rect 18478 20479 18536 20485
rect 13504 20411 13516 20457
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 15861 20451 15919 20457
rect 15861 20417 15873 20451
rect 15907 20448 15919 20451
rect 16758 20448 16764 20460
rect 15907 20420 16764 20448
rect 15907 20417 15919 20420
rect 15861 20411 15919 20417
rect 13504 20408 13510 20411
rect 16758 20408 16764 20420
rect 16816 20408 16822 20460
rect 17310 20408 17316 20460
rect 17368 20448 17374 20460
rect 17874 20451 17932 20457
rect 17874 20448 17886 20451
rect 17368 20420 17886 20448
rect 17368 20408 17374 20420
rect 17874 20417 17886 20420
rect 17920 20417 17932 20451
rect 17874 20411 17932 20417
rect 6270 20340 6276 20392
rect 6328 20380 6334 20392
rect 6733 20383 6791 20389
rect 6733 20380 6745 20383
rect 6328 20352 6745 20380
rect 6328 20340 6334 20352
rect 6733 20349 6745 20352
rect 6779 20349 6791 20383
rect 6733 20343 6791 20349
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 8386 20380 8392 20392
rect 7055 20352 8392 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 3878 20204 3884 20256
rect 3936 20204 3942 20256
rect 6641 20247 6699 20253
rect 6641 20213 6653 20247
rect 6687 20244 6699 20247
rect 6748 20244 6776 20343
rect 8386 20340 8392 20352
rect 8444 20340 8450 20392
rect 10042 20340 10048 20392
rect 10100 20340 10106 20392
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20349 10379 20383
rect 10321 20343 10379 20349
rect 7006 20244 7012 20256
rect 6687 20216 7012 20244
rect 6687 20213 6699 20216
rect 6641 20207 6699 20213
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 8570 20204 8576 20256
rect 8628 20204 8634 20256
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 10336 20244 10364 20343
rect 16114 20340 16120 20392
rect 16172 20340 16178 20392
rect 18141 20383 18199 20389
rect 18141 20349 18153 20383
rect 18187 20380 18199 20383
rect 18233 20383 18291 20389
rect 18233 20380 18245 20383
rect 18187 20352 18245 20380
rect 18187 20349 18199 20352
rect 18141 20343 18199 20349
rect 18233 20349 18245 20352
rect 18279 20349 18291 20383
rect 18233 20343 18291 20349
rect 9732 20216 10364 20244
rect 9732 20204 9738 20216
rect 12342 20204 12348 20256
rect 12400 20204 12406 20256
rect 14734 20204 14740 20256
rect 14792 20204 14798 20256
rect 15378 20204 15384 20256
rect 15436 20244 15442 20256
rect 16132 20244 16160 20340
rect 15436 20216 16160 20244
rect 16761 20247 16819 20253
rect 15436 20204 15442 20216
rect 16761 20213 16773 20247
rect 16807 20244 16819 20247
rect 17126 20244 17132 20256
rect 16807 20216 17132 20244
rect 16807 20213 16819 20216
rect 16761 20207 16819 20213
rect 17126 20204 17132 20216
rect 17184 20204 17190 20256
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 18156 20244 18184 20343
rect 18012 20216 18184 20244
rect 19613 20247 19671 20253
rect 18012 20204 18018 20216
rect 19613 20213 19625 20247
rect 19659 20244 19671 20247
rect 19794 20244 19800 20256
rect 19659 20216 19800 20244
rect 19659 20213 19671 20216
rect 19613 20207 19671 20213
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 1104 20154 20792 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 10214 20154
rect 10266 20102 10278 20154
rect 10330 20102 10342 20154
rect 10394 20102 10406 20154
rect 10458 20102 10470 20154
rect 10522 20102 16214 20154
rect 16266 20102 16278 20154
rect 16330 20102 16342 20154
rect 16394 20102 16406 20154
rect 16458 20102 16470 20154
rect 16522 20102 20792 20154
rect 1104 20080 20792 20102
rect 3878 20000 3884 20052
rect 3936 20000 3942 20052
rect 5997 20043 6055 20049
rect 5997 20009 6009 20043
rect 6043 20040 6055 20043
rect 6270 20040 6276 20052
rect 6043 20012 6276 20040
rect 6043 20009 6055 20012
rect 5997 20003 6055 20009
rect 6270 20000 6276 20012
rect 6328 20000 6334 20052
rect 8386 20000 8392 20052
rect 8444 20000 8450 20052
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 10229 20043 10287 20049
rect 10229 20040 10241 20043
rect 10100 20012 10241 20040
rect 10100 20000 10106 20012
rect 10229 20009 10241 20012
rect 10275 20009 10287 20043
rect 10229 20003 10287 20009
rect 13446 20000 13452 20052
rect 13504 20040 13510 20052
rect 13541 20043 13599 20049
rect 13541 20040 13553 20043
rect 13504 20012 13553 20040
rect 13504 20000 13510 20012
rect 13541 20009 13553 20012
rect 13587 20040 13599 20043
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 13587 20012 14105 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 14093 20003 14151 20009
rect 14734 20000 14740 20052
rect 14792 20000 14798 20052
rect 3896 19845 3924 20000
rect 6365 19975 6423 19981
rect 6365 19941 6377 19975
rect 6411 19972 6423 19975
rect 6411 19944 6500 19972
rect 6411 19941 6423 19944
rect 6365 19935 6423 19941
rect 6472 19913 6500 19944
rect 6457 19907 6515 19913
rect 6457 19873 6469 19907
rect 6503 19873 6515 19907
rect 9398 19904 9404 19916
rect 6457 19867 6515 19873
rect 6932 19876 7420 19904
rect 6932 19848 6960 19876
rect 3881 19839 3939 19845
rect 3881 19805 3893 19839
rect 3927 19805 3939 19839
rect 3881 19799 3939 19805
rect 6089 19839 6147 19845
rect 6089 19805 6101 19839
rect 6135 19805 6147 19839
rect 6089 19799 6147 19805
rect 6104 19712 6132 19799
rect 6914 19796 6920 19848
rect 6972 19796 6978 19848
rect 7392 19845 7420 19876
rect 8496 19876 9404 19904
rect 8496 19845 8524 19876
rect 9398 19864 9404 19876
rect 9456 19904 9462 19916
rect 9769 19907 9827 19913
rect 9769 19904 9781 19907
rect 9456 19876 9781 19904
rect 9456 19864 9462 19876
rect 9769 19873 9781 19876
rect 9815 19873 9827 19907
rect 14752 19904 14780 20000
rect 14752 19876 15516 19904
rect 9769 19867 9827 19873
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 7193 19839 7251 19845
rect 7193 19836 7205 19839
rect 7147 19808 7205 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 7193 19805 7205 19808
rect 7239 19805 7251 19839
rect 7193 19799 7251 19805
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19805 7435 19839
rect 7377 19799 7435 19805
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19805 8539 19839
rect 8481 19799 8539 19805
rect 8570 19796 8576 19848
rect 8628 19836 8634 19848
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 8628 19808 8953 19836
rect 8628 19796 8634 19808
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 8941 19799 8999 19805
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19836 9643 19839
rect 9861 19839 9919 19845
rect 9861 19836 9873 19839
rect 9631 19808 9873 19836
rect 9631 19805 9643 19808
rect 9585 19799 9643 19805
rect 9861 19805 9873 19808
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 11514 19796 11520 19848
rect 11572 19836 11578 19848
rect 12434 19845 12440 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11572 19808 12173 19836
rect 11572 19796 11578 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12428 19799 12440 19845
rect 12492 19836 12498 19848
rect 13630 19836 13636 19848
rect 12492 19808 13636 19836
rect 12434 19796 12440 19799
rect 12492 19796 12498 19808
rect 13630 19796 13636 19808
rect 13688 19836 13694 19848
rect 14093 19839 14151 19845
rect 14093 19836 14105 19839
rect 13688 19808 14105 19836
rect 13688 19796 13694 19808
rect 14093 19805 14105 19808
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 14182 19796 14188 19848
rect 14240 19796 14246 19848
rect 15286 19796 15292 19848
rect 15344 19836 15350 19848
rect 15381 19839 15439 19845
rect 15381 19836 15393 19839
rect 15344 19808 15393 19836
rect 15344 19796 15350 19808
rect 15381 19805 15393 19808
rect 15427 19805 15439 19839
rect 15488 19836 15516 19876
rect 16684 19876 17448 19904
rect 15637 19839 15695 19845
rect 15637 19836 15649 19839
rect 15488 19808 15649 19836
rect 15381 19799 15439 19805
rect 15637 19805 15649 19808
rect 15683 19836 15695 19839
rect 16684 19836 16712 19876
rect 17221 19839 17279 19845
rect 17221 19836 17233 19839
rect 15683 19808 16712 19836
rect 16776 19808 17233 19836
rect 15683 19805 15695 19808
rect 15637 19799 15695 19805
rect 6362 19728 6368 19780
rect 6420 19728 6426 19780
rect 3510 19660 3516 19712
rect 3568 19700 3574 19712
rect 3881 19703 3939 19709
rect 3881 19700 3893 19703
rect 3568 19672 3893 19700
rect 3568 19660 3574 19672
rect 3881 19669 3893 19672
rect 3927 19669 3939 19703
rect 3881 19663 3939 19669
rect 6086 19660 6092 19712
rect 6144 19660 6150 19712
rect 6178 19660 6184 19712
rect 6236 19660 6242 19712
rect 7285 19703 7343 19709
rect 7285 19669 7297 19703
rect 7331 19700 7343 19703
rect 7558 19700 7564 19712
rect 7331 19672 7564 19700
rect 7331 19669 7343 19672
rect 7285 19663 7343 19669
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 14458 19660 14464 19712
rect 14516 19660 14522 19712
rect 16776 19709 16804 19808
rect 17221 19805 17233 19808
rect 17267 19836 17279 19839
rect 17310 19836 17316 19848
rect 17267 19808 17316 19836
rect 17267 19805 17279 19808
rect 17221 19799 17279 19805
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 16945 19771 17003 19777
rect 16945 19737 16957 19771
rect 16991 19768 17003 19771
rect 17034 19768 17040 19780
rect 16991 19740 17040 19768
rect 16991 19737 17003 19740
rect 16945 19731 17003 19737
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 17420 19712 17448 19876
rect 17954 19796 17960 19848
rect 18012 19836 18018 19848
rect 19061 19839 19119 19845
rect 19061 19836 19073 19839
rect 18012 19808 19073 19836
rect 18012 19796 18018 19808
rect 19061 19805 19073 19808
rect 19107 19805 19119 19839
rect 19061 19799 19119 19805
rect 18816 19771 18874 19777
rect 18816 19737 18828 19771
rect 18862 19768 18874 19771
rect 19794 19768 19800 19780
rect 18862 19740 19800 19768
rect 18862 19737 18874 19740
rect 18816 19731 18874 19737
rect 19794 19728 19800 19740
rect 19852 19728 19858 19780
rect 16761 19703 16819 19709
rect 16761 19669 16773 19703
rect 16807 19669 16819 19703
rect 16761 19663 16819 19669
rect 17126 19660 17132 19712
rect 17184 19660 17190 19712
rect 17313 19703 17371 19709
rect 17313 19669 17325 19703
rect 17359 19700 17371 19703
rect 17402 19700 17408 19712
rect 17359 19672 17408 19700
rect 17359 19669 17371 19672
rect 17313 19663 17371 19669
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 17494 19660 17500 19712
rect 17552 19660 17558 19712
rect 17678 19660 17684 19712
rect 17736 19660 17742 19712
rect 1104 19610 20792 19632
rect 1104 19558 7214 19610
rect 7266 19558 7278 19610
rect 7330 19558 7342 19610
rect 7394 19558 7406 19610
rect 7458 19558 7470 19610
rect 7522 19558 13214 19610
rect 13266 19558 13278 19610
rect 13330 19558 13342 19610
rect 13394 19558 13406 19610
rect 13458 19558 13470 19610
rect 13522 19558 19214 19610
rect 19266 19558 19278 19610
rect 19330 19558 19342 19610
rect 19394 19558 19406 19610
rect 19458 19558 19470 19610
rect 19522 19558 20792 19610
rect 1104 19536 20792 19558
rect 4617 19499 4675 19505
rect 4617 19465 4629 19499
rect 4663 19496 4675 19499
rect 6270 19496 6276 19508
rect 4663 19468 6276 19496
rect 4663 19465 4675 19468
rect 4617 19459 4675 19465
rect 4249 19431 4307 19437
rect 4249 19428 4261 19431
rect 3160 19400 4261 19428
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19360 2559 19363
rect 2774 19360 2780 19372
rect 2547 19332 2780 19360
rect 2547 19329 2559 19332
rect 2501 19323 2559 19329
rect 2774 19320 2780 19332
rect 2832 19320 2838 19372
rect 3160 19369 3188 19400
rect 4249 19397 4261 19400
rect 4295 19397 4307 19431
rect 4249 19391 4307 19397
rect 3145 19363 3203 19369
rect 3145 19329 3157 19363
rect 3191 19329 3203 19363
rect 3145 19323 3203 19329
rect 3237 19363 3295 19369
rect 3237 19329 3249 19363
rect 3283 19360 3295 19363
rect 3510 19360 3516 19372
rect 3283 19332 3516 19360
rect 3283 19329 3295 19332
rect 3237 19323 3295 19329
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 4724 19369 4752 19468
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 6362 19456 6368 19508
rect 6420 19496 6426 19508
rect 6457 19499 6515 19505
rect 6457 19496 6469 19499
rect 6420 19468 6469 19496
rect 6420 19456 6426 19468
rect 6457 19465 6469 19468
rect 6503 19465 6515 19499
rect 6457 19459 6515 19465
rect 8570 19456 8576 19508
rect 8628 19496 8634 19508
rect 10137 19499 10195 19505
rect 10137 19496 10149 19499
rect 8628 19468 10149 19496
rect 8628 19456 8634 19468
rect 10137 19465 10149 19468
rect 10183 19465 10195 19499
rect 10137 19459 10195 19465
rect 11514 19456 11520 19508
rect 11572 19496 11578 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 11572 19468 11805 19496
rect 11572 19456 11578 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 11793 19459 11851 19465
rect 13078 19456 13084 19508
rect 13136 19496 13142 19508
rect 13357 19499 13415 19505
rect 13357 19496 13369 19499
rect 13136 19468 13369 19496
rect 13136 19456 13142 19468
rect 13357 19465 13369 19468
rect 13403 19465 13415 19499
rect 14182 19496 14188 19508
rect 13357 19459 13415 19465
rect 13464 19468 14188 19496
rect 7558 19388 7564 19440
rect 7616 19437 7622 19440
rect 7616 19428 7628 19437
rect 9309 19431 9367 19437
rect 9309 19428 9321 19431
rect 7616 19400 7661 19428
rect 9232 19400 9321 19428
rect 7616 19391 7628 19400
rect 7616 19388 7622 19391
rect 4982 19369 4988 19372
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19329 4031 19363
rect 3973 19323 4031 19329
rect 4709 19363 4767 19369
rect 4709 19329 4721 19363
rect 4755 19329 4767 19363
rect 4709 19323 4767 19329
rect 4976 19323 4988 19369
rect 3881 19295 3939 19301
rect 3881 19261 3893 19295
rect 3927 19292 3939 19295
rect 3988 19292 4016 19323
rect 4982 19320 4988 19323
rect 5040 19320 5046 19372
rect 9033 19363 9091 19369
rect 9033 19329 9045 19363
rect 9079 19360 9091 19363
rect 9122 19360 9128 19372
rect 9079 19332 9128 19360
rect 9079 19329 9091 19332
rect 9033 19323 9091 19329
rect 9122 19320 9128 19332
rect 9180 19320 9186 19372
rect 9232 19369 9260 19400
rect 9309 19397 9321 19400
rect 9355 19397 9367 19431
rect 9309 19391 9367 19397
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 13464 19428 13492 19468
rect 12400 19400 13492 19428
rect 13525 19431 13583 19437
rect 12400 19388 12406 19400
rect 13525 19397 13537 19431
rect 13571 19428 13583 19431
rect 13630 19428 13636 19440
rect 13571 19400 13636 19428
rect 13571 19397 13583 19400
rect 13525 19391 13583 19397
rect 13630 19388 13636 19400
rect 13688 19388 13694 19440
rect 13725 19431 13783 19437
rect 13725 19397 13737 19431
rect 13771 19428 13783 19431
rect 13832 19428 13860 19468
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 16117 19499 16175 19505
rect 16117 19465 16129 19499
rect 16163 19496 16175 19499
rect 16942 19496 16948 19508
rect 16163 19468 16948 19496
rect 16163 19465 16175 19468
rect 16117 19459 16175 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 16574 19428 16580 19440
rect 13771 19400 13860 19428
rect 15304 19400 16580 19428
rect 13771 19397 13783 19400
rect 13725 19391 13783 19397
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19329 9275 19363
rect 9217 19323 9275 19329
rect 9582 19320 9588 19372
rect 9640 19360 9646 19372
rect 10045 19363 10103 19369
rect 10045 19360 10057 19363
rect 9640 19332 10057 19360
rect 9640 19320 9646 19332
rect 10045 19329 10057 19332
rect 10091 19329 10103 19363
rect 10045 19323 10103 19329
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10505 19363 10563 19369
rect 10505 19360 10517 19363
rect 10367 19332 10517 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10505 19329 10517 19332
rect 10551 19329 10563 19363
rect 10505 19323 10563 19329
rect 13265 19363 13323 19369
rect 13265 19329 13277 19363
rect 13311 19360 13323 19363
rect 15304 19360 15332 19400
rect 16574 19388 16580 19400
rect 16632 19428 16638 19440
rect 16669 19431 16727 19437
rect 16669 19428 16681 19431
rect 16632 19400 16681 19428
rect 16632 19388 16638 19400
rect 16669 19397 16681 19400
rect 16715 19397 16727 19431
rect 16669 19391 16727 19397
rect 13311 19332 15332 19360
rect 16485 19363 16543 19369
rect 13311 19329 13323 19332
rect 13265 19323 13323 19329
rect 16485 19329 16497 19363
rect 16531 19360 16543 19363
rect 18046 19360 18052 19372
rect 16531 19332 18052 19360
rect 16531 19329 16543 19332
rect 16485 19323 16543 19329
rect 18046 19320 18052 19332
rect 18104 19320 18110 19372
rect 18782 19369 18788 19372
rect 18776 19323 18788 19369
rect 18782 19320 18788 19323
rect 18840 19320 18846 19372
rect 3927 19264 4016 19292
rect 3927 19261 3939 19264
rect 3881 19255 3939 19261
rect 7834 19252 7840 19304
rect 7892 19292 7898 19304
rect 9306 19292 9312 19304
rect 7892 19264 9312 19292
rect 7892 19252 7898 19264
rect 9306 19252 9312 19264
rect 9364 19292 9370 19304
rect 9674 19292 9680 19304
rect 9364 19264 9680 19292
rect 9364 19252 9370 19264
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19261 9919 19295
rect 9861 19255 9919 19261
rect 6089 19227 6147 19233
rect 6089 19193 6101 19227
rect 6135 19224 6147 19227
rect 6178 19224 6184 19236
rect 6135 19196 6184 19224
rect 6135 19193 6147 19196
rect 6089 19187 6147 19193
rect 6178 19184 6184 19196
rect 6236 19184 6242 19236
rect 8754 19184 8760 19236
rect 8812 19224 8818 19236
rect 9214 19224 9220 19236
rect 8812 19196 9220 19224
rect 8812 19184 8818 19196
rect 9214 19184 9220 19196
rect 9272 19224 9278 19236
rect 9876 19224 9904 19255
rect 11146 19252 11152 19304
rect 11204 19252 11210 19304
rect 16393 19295 16451 19301
rect 16393 19261 16405 19295
rect 16439 19292 16451 19295
rect 16666 19292 16672 19304
rect 16439 19264 16672 19292
rect 16439 19261 16451 19264
rect 16393 19255 16451 19261
rect 16666 19252 16672 19264
rect 16724 19252 16730 19304
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 17972 19264 18521 19292
rect 9272 19196 9904 19224
rect 9272 19184 9278 19196
rect 17972 19168 18000 19264
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 18509 19255 18567 19261
rect 9030 19116 9036 19168
rect 9088 19116 9094 19168
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 10321 19159 10379 19165
rect 10321 19156 10333 19159
rect 10100 19128 10333 19156
rect 10100 19116 10106 19128
rect 10321 19125 10333 19128
rect 10367 19125 10379 19159
rect 10321 19119 10379 19125
rect 13538 19116 13544 19168
rect 13596 19116 13602 19168
rect 16485 19159 16543 19165
rect 16485 19125 16497 19159
rect 16531 19156 16543 19159
rect 16850 19156 16856 19168
rect 16531 19128 16856 19156
rect 16531 19125 16543 19128
rect 16485 19119 16543 19125
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 17954 19116 17960 19168
rect 18012 19116 18018 19168
rect 19886 19116 19892 19168
rect 19944 19116 19950 19168
rect 1104 19066 20792 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 10214 19066
rect 10266 19014 10278 19066
rect 10330 19014 10342 19066
rect 10394 19014 10406 19066
rect 10458 19014 10470 19066
rect 10522 19014 16214 19066
rect 16266 19014 16278 19066
rect 16330 19014 16342 19066
rect 16394 19014 16406 19066
rect 16458 19014 16470 19066
rect 16522 19014 20792 19066
rect 1104 18992 20792 19014
rect 4982 18912 4988 18964
rect 5040 18952 5046 18964
rect 5077 18955 5135 18961
rect 5077 18952 5089 18955
rect 5040 18924 5089 18952
rect 5040 18912 5046 18924
rect 5077 18921 5089 18924
rect 5123 18921 5135 18955
rect 5077 18915 5135 18921
rect 6362 18912 6368 18964
rect 6420 18952 6426 18964
rect 6641 18955 6699 18961
rect 6641 18952 6653 18955
rect 6420 18924 6653 18952
rect 6420 18912 6426 18924
rect 6641 18921 6653 18924
rect 6687 18921 6699 18955
rect 6641 18915 6699 18921
rect 6825 18955 6883 18961
rect 6825 18921 6837 18955
rect 6871 18952 6883 18955
rect 6914 18952 6920 18964
rect 6871 18924 6920 18952
rect 6871 18921 6883 18924
rect 6825 18915 6883 18921
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 8754 18912 8760 18964
rect 8812 18912 8818 18964
rect 9122 18912 9128 18964
rect 9180 18912 9186 18964
rect 9217 18955 9275 18961
rect 9217 18921 9229 18955
rect 9263 18952 9275 18955
rect 9582 18952 9588 18964
rect 9263 18924 9588 18952
rect 9263 18921 9275 18924
rect 9217 18915 9275 18921
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11241 18955 11299 18961
rect 11241 18952 11253 18955
rect 11204 18924 11253 18952
rect 11204 18912 11210 18924
rect 11241 18921 11253 18924
rect 11287 18921 11299 18955
rect 11241 18915 11299 18921
rect 16669 18955 16727 18961
rect 16669 18921 16681 18955
rect 16715 18952 16727 18955
rect 16758 18952 16764 18964
rect 16715 18924 16764 18952
rect 16715 18921 16727 18924
rect 16669 18915 16727 18921
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 16850 18912 16856 18964
rect 16908 18912 16914 18964
rect 17126 18912 17132 18964
rect 17184 18912 17190 18964
rect 18782 18912 18788 18964
rect 18840 18952 18846 18964
rect 18969 18955 19027 18961
rect 18969 18952 18981 18955
rect 18840 18924 18981 18952
rect 18840 18912 18846 18924
rect 18969 18921 18981 18924
rect 19015 18921 19027 18955
rect 18969 18915 19027 18921
rect 2777 18887 2835 18893
rect 2777 18853 2789 18887
rect 2823 18853 2835 18887
rect 9140 18884 9168 18912
rect 9401 18887 9459 18893
rect 9401 18884 9413 18887
rect 9140 18856 9413 18884
rect 2777 18847 2835 18853
rect 9401 18853 9413 18856
rect 9447 18884 9459 18887
rect 9490 18884 9496 18896
rect 9447 18856 9496 18884
rect 9447 18853 9459 18856
rect 9401 18847 9459 18853
rect 2792 18816 2820 18847
rect 9490 18844 9496 18856
rect 9548 18844 9554 18896
rect 2700 18788 2820 18816
rect 5721 18819 5779 18825
rect 2700 18757 2728 18788
rect 5721 18785 5733 18819
rect 5767 18816 5779 18819
rect 5813 18819 5871 18825
rect 5813 18816 5825 18819
rect 5767 18788 5825 18816
rect 5767 18785 5779 18788
rect 5721 18779 5779 18785
rect 5813 18785 5825 18788
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 6086 18776 6092 18828
rect 6144 18816 6150 18828
rect 6144 18788 6592 18816
rect 6144 18776 6150 18788
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18717 2743 18751
rect 2685 18711 2743 18717
rect 2774 18708 2780 18760
rect 2832 18708 2838 18760
rect 6178 18708 6184 18760
rect 6236 18708 6242 18760
rect 6196 18680 6224 18708
rect 6457 18683 6515 18689
rect 6457 18680 6469 18683
rect 6196 18652 6469 18680
rect 6457 18649 6469 18652
rect 6503 18649 6515 18683
rect 6564 18680 6592 18788
rect 7006 18776 7012 18828
rect 7064 18816 7070 18828
rect 7834 18816 7840 18828
rect 7064 18788 7840 18816
rect 7064 18776 7070 18788
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 8846 18816 8852 18828
rect 8404 18788 8852 18816
rect 8294 18708 8300 18760
rect 8352 18748 8358 18760
rect 8404 18748 8432 18788
rect 8846 18776 8852 18788
rect 8904 18816 8910 18828
rect 8904 18788 10916 18816
rect 8904 18776 8910 18788
rect 8352 18734 8432 18748
rect 8352 18720 8418 18734
rect 8352 18708 8358 18720
rect 9306 18708 9312 18760
rect 9364 18748 9370 18760
rect 9493 18751 9551 18757
rect 9493 18748 9505 18751
rect 9364 18720 9505 18748
rect 9364 18708 9370 18720
rect 9493 18717 9505 18720
rect 9539 18717 9551 18751
rect 10888 18734 10916 18788
rect 9493 18711 9551 18717
rect 6657 18683 6715 18689
rect 6657 18680 6669 18683
rect 6564 18652 6669 18680
rect 6457 18643 6515 18649
rect 6657 18649 6669 18652
rect 6703 18649 6715 18683
rect 6657 18643 6715 18649
rect 7285 18683 7343 18689
rect 7285 18649 7297 18683
rect 7331 18680 7343 18683
rect 7558 18680 7564 18692
rect 7331 18652 7564 18680
rect 7331 18649 7343 18652
rect 7285 18643 7343 18649
rect 7558 18640 7564 18652
rect 7616 18640 7622 18692
rect 8570 18640 8576 18692
rect 8628 18680 8634 18692
rect 9033 18683 9091 18689
rect 9033 18680 9045 18683
rect 8628 18652 9045 18680
rect 8628 18640 8634 18652
rect 9033 18649 9045 18652
rect 9079 18680 9091 18683
rect 9122 18680 9128 18692
rect 9079 18652 9128 18680
rect 9079 18649 9091 18652
rect 9033 18643 9091 18649
rect 9122 18640 9128 18652
rect 9180 18640 9186 18692
rect 9766 18640 9772 18692
rect 9824 18640 9830 18692
rect 2038 18572 2044 18624
rect 2096 18572 2102 18624
rect 9243 18615 9301 18621
rect 9243 18581 9255 18615
rect 9289 18612 9301 18615
rect 9398 18612 9404 18624
rect 9289 18584 9404 18612
rect 9289 18581 9301 18584
rect 9243 18575 9301 18581
rect 9398 18572 9404 18584
rect 9456 18612 9462 18624
rect 11164 18612 11192 18912
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11609 18819 11667 18825
rect 11609 18816 11621 18819
rect 11572 18788 11621 18816
rect 11572 18776 11578 18788
rect 11609 18785 11621 18788
rect 11655 18785 11667 18819
rect 11609 18779 11667 18785
rect 17589 18819 17647 18825
rect 17589 18785 17601 18819
rect 17635 18785 17647 18819
rect 17589 18779 17647 18785
rect 11876 18751 11934 18757
rect 11876 18717 11888 18751
rect 11922 18748 11934 18751
rect 12342 18748 12348 18760
rect 11922 18720 12348 18748
rect 11922 18717 11934 18720
rect 11876 18711 11934 18717
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 15286 18708 15292 18760
rect 15344 18708 15350 18760
rect 15556 18751 15614 18757
rect 15556 18717 15568 18751
rect 15602 18717 15614 18751
rect 15556 18711 15614 18717
rect 9456 18584 11192 18612
rect 9456 18572 9462 18584
rect 12986 18572 12992 18624
rect 13044 18572 13050 18624
rect 15304 18612 15332 18708
rect 15470 18640 15476 18692
rect 15528 18680 15534 18692
rect 15580 18680 15608 18711
rect 17034 18708 17040 18760
rect 17092 18708 17098 18760
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 17218 18748 17224 18760
rect 17175 18720 17224 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18748 17371 18751
rect 17402 18748 17408 18760
rect 17359 18720 17408 18748
rect 17359 18717 17371 18720
rect 17313 18711 17371 18717
rect 17402 18708 17408 18720
rect 17460 18708 17466 18760
rect 17604 18680 17632 18779
rect 17678 18708 17684 18760
rect 17736 18748 17742 18760
rect 17845 18751 17903 18757
rect 17845 18748 17857 18751
rect 17736 18720 17857 18748
rect 17736 18708 17742 18720
rect 17845 18717 17857 18720
rect 17891 18748 17903 18751
rect 18984 18748 19012 18915
rect 19886 18844 19892 18896
rect 19944 18884 19950 18896
rect 20257 18887 20315 18893
rect 20257 18884 20269 18887
rect 19944 18856 20269 18884
rect 19944 18844 19950 18856
rect 20257 18853 20269 18856
rect 20303 18853 20315 18887
rect 20257 18847 20315 18853
rect 19610 18748 19616 18760
rect 17891 18720 18828 18748
rect 18984 18720 19616 18748
rect 17891 18717 17903 18720
rect 17845 18711 17903 18717
rect 17954 18680 17960 18692
rect 15528 18652 15608 18680
rect 16132 18652 17960 18680
rect 15528 18640 15534 18652
rect 16132 18624 16160 18652
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 18800 18680 18828 18720
rect 19610 18708 19616 18720
rect 19668 18748 19674 18760
rect 20073 18751 20131 18757
rect 20073 18748 20085 18751
rect 19668 18720 20085 18748
rect 19668 18708 19674 18720
rect 20073 18717 20085 18720
rect 20119 18717 20131 18751
rect 20073 18711 20131 18717
rect 19978 18680 19984 18692
rect 18800 18652 19984 18680
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 16114 18612 16120 18624
rect 15304 18584 16120 18612
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 19702 18572 19708 18624
rect 19760 18572 19766 18624
rect 19794 18572 19800 18624
rect 19852 18612 19858 18624
rect 19889 18615 19947 18621
rect 19889 18612 19901 18615
rect 19852 18584 19901 18612
rect 19852 18572 19858 18584
rect 19889 18581 19901 18584
rect 19935 18581 19947 18615
rect 19889 18575 19947 18581
rect 1104 18522 20792 18544
rect 1104 18470 7214 18522
rect 7266 18470 7278 18522
rect 7330 18470 7342 18522
rect 7394 18470 7406 18522
rect 7458 18470 7470 18522
rect 7522 18470 13214 18522
rect 13266 18470 13278 18522
rect 13330 18470 13342 18522
rect 13394 18470 13406 18522
rect 13458 18470 13470 18522
rect 13522 18470 19214 18522
rect 19266 18470 19278 18522
rect 19330 18470 19342 18522
rect 19394 18470 19406 18522
rect 19458 18470 19470 18522
rect 19522 18470 20792 18522
rect 1104 18448 20792 18470
rect 2038 18368 2044 18420
rect 2096 18368 2102 18420
rect 6917 18411 6975 18417
rect 6917 18377 6929 18411
rect 6963 18408 6975 18411
rect 7006 18408 7012 18420
rect 6963 18380 7012 18408
rect 6963 18377 6975 18380
rect 6917 18371 6975 18377
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 8849 18411 8907 18417
rect 8849 18408 8861 18411
rect 7616 18380 8861 18408
rect 7616 18368 7622 18380
rect 8849 18377 8861 18380
rect 8895 18377 8907 18411
rect 8849 18371 8907 18377
rect 9030 18368 9036 18420
rect 9088 18368 9094 18420
rect 9214 18368 9220 18420
rect 9272 18368 9278 18420
rect 9309 18411 9367 18417
rect 9309 18377 9321 18411
rect 9355 18408 9367 18411
rect 9398 18408 9404 18420
rect 9355 18380 9404 18408
rect 9355 18377 9367 18380
rect 9309 18371 9367 18377
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 9766 18368 9772 18420
rect 9824 18368 9830 18420
rect 15381 18411 15439 18417
rect 15381 18377 15393 18411
rect 15427 18377 15439 18411
rect 15381 18371 15439 18377
rect 2056 18272 2084 18368
rect 9048 18340 9076 18368
rect 8772 18312 9076 18340
rect 8772 18281 8800 18312
rect 9122 18300 9128 18352
rect 9180 18340 9186 18352
rect 9585 18343 9643 18349
rect 9585 18340 9597 18343
rect 9180 18312 9597 18340
rect 9180 18300 9186 18312
rect 9585 18309 9597 18312
rect 9631 18309 9643 18343
rect 9585 18303 9643 18309
rect 12986 18300 12992 18352
rect 13044 18340 13050 18352
rect 13446 18340 13452 18352
rect 13044 18312 13452 18340
rect 13044 18300 13050 18312
rect 13446 18300 13452 18312
rect 13504 18340 13510 18352
rect 14274 18349 14280 18352
rect 13642 18343 13700 18349
rect 13642 18340 13654 18343
rect 13504 18312 13654 18340
rect 13504 18300 13510 18312
rect 13642 18309 13654 18312
rect 13688 18309 13700 18343
rect 14268 18340 14280 18349
rect 14235 18312 14280 18340
rect 13642 18303 13700 18309
rect 14268 18303 14280 18312
rect 14274 18300 14280 18303
rect 14332 18300 14338 18352
rect 15396 18340 15424 18371
rect 16666 18368 16672 18420
rect 16724 18368 16730 18420
rect 17681 18411 17739 18417
rect 17681 18408 17693 18411
rect 17236 18380 17693 18408
rect 15838 18340 15844 18352
rect 15396 18312 15844 18340
rect 15838 18300 15844 18312
rect 15896 18340 15902 18352
rect 17236 18349 17264 18380
rect 17681 18377 17693 18380
rect 17727 18377 17739 18411
rect 19702 18408 19708 18420
rect 17681 18371 17739 18377
rect 17788 18380 19708 18408
rect 17221 18343 17279 18349
rect 15896 18312 17080 18340
rect 15896 18300 15902 18312
rect 2133 18275 2191 18281
rect 2133 18272 2145 18275
rect 2056 18244 2145 18272
rect 2133 18241 2145 18244
rect 2179 18241 2191 18275
rect 2133 18235 2191 18241
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18241 8815 18275
rect 8757 18235 8815 18241
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18272 8999 18275
rect 9033 18275 9091 18281
rect 9033 18272 9045 18275
rect 8987 18244 9045 18272
rect 8987 18241 8999 18244
rect 8941 18235 8999 18241
rect 9033 18241 9045 18244
rect 9079 18241 9091 18275
rect 9033 18235 9091 18241
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18241 9459 18275
rect 9401 18235 9459 18241
rect 9048 18136 9076 18235
rect 9416 18204 9444 18235
rect 9490 18232 9496 18284
rect 9548 18272 9554 18284
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9548 18244 9689 18272
rect 9548 18232 9554 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18272 9919 18275
rect 10042 18272 10048 18284
rect 9907 18244 10048 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 13909 18275 13967 18281
rect 13909 18272 13921 18275
rect 13872 18244 13921 18272
rect 13872 18232 13878 18244
rect 13909 18241 13921 18244
rect 13955 18272 13967 18275
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13955 18244 14013 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 17052 18281 17080 18312
rect 17221 18309 17233 18343
rect 17267 18309 17279 18343
rect 17221 18303 17279 18309
rect 17437 18343 17495 18349
rect 17437 18309 17449 18343
rect 17483 18340 17495 18343
rect 17788 18340 17816 18380
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 17483 18312 17816 18340
rect 17849 18343 17907 18349
rect 17483 18309 17495 18312
rect 17437 18303 17495 18309
rect 17849 18309 17861 18343
rect 17895 18309 17907 18343
rect 17849 18303 17907 18309
rect 18049 18343 18107 18349
rect 18049 18309 18061 18343
rect 18095 18309 18107 18343
rect 18049 18303 18107 18309
rect 18868 18343 18926 18349
rect 18868 18309 18880 18343
rect 18914 18340 18926 18343
rect 19426 18340 19432 18352
rect 18914 18312 19432 18340
rect 18914 18309 18926 18312
rect 18868 18303 18926 18309
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16816 18244 16865 18272
rect 16816 18232 16822 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17037 18275 17095 18281
rect 17037 18241 17049 18275
rect 17083 18272 17095 18275
rect 17871 18272 17899 18303
rect 17083 18244 17899 18272
rect 17083 18241 17095 18244
rect 17037 18235 17095 18241
rect 9582 18204 9588 18216
rect 9416 18176 9588 18204
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 16868 18204 16896 18235
rect 18064 18204 18092 18303
rect 19426 18300 19432 18312
rect 19484 18340 19490 18352
rect 19886 18340 19892 18352
rect 19484 18312 19892 18340
rect 19484 18300 19490 18312
rect 19886 18300 19892 18312
rect 19944 18300 19950 18352
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 16868 18176 18092 18204
rect 9490 18136 9496 18148
rect 9048 18108 9496 18136
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 17328 18108 17908 18136
rect 2130 18028 2136 18080
rect 2188 18028 2194 18080
rect 9306 18028 9312 18080
rect 9364 18068 9370 18080
rect 10229 18071 10287 18077
rect 10229 18068 10241 18071
rect 9364 18040 10241 18068
rect 9364 18028 9370 18040
rect 10229 18037 10241 18040
rect 10275 18037 10287 18071
rect 10229 18031 10287 18037
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 13170 18068 13176 18080
rect 12584 18040 13176 18068
rect 12584 18028 12590 18040
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 15528 18040 16865 18068
rect 15528 18028 15534 18040
rect 16853 18037 16865 18040
rect 16899 18068 16911 18071
rect 17328 18068 17356 18108
rect 16899 18040 17356 18068
rect 17405 18071 17463 18077
rect 16899 18037 16911 18040
rect 16853 18031 16911 18037
rect 17405 18037 17417 18071
rect 17451 18068 17463 18071
rect 17494 18068 17500 18080
rect 17451 18040 17500 18068
rect 17451 18037 17463 18040
rect 17405 18031 17463 18037
rect 17494 18028 17500 18040
rect 17552 18028 17558 18080
rect 17586 18028 17592 18080
rect 17644 18028 17650 18080
rect 17880 18077 17908 18108
rect 17954 18096 17960 18148
rect 18012 18136 18018 18148
rect 18616 18136 18644 18235
rect 18012 18108 18644 18136
rect 18012 18096 18018 18108
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18037 17923 18071
rect 17865 18031 17923 18037
rect 19702 18028 19708 18080
rect 19760 18068 19766 18080
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 19760 18040 19993 18068
rect 19760 18028 19766 18040
rect 19981 18037 19993 18040
rect 20027 18037 20039 18071
rect 19981 18031 20039 18037
rect 1104 17978 20792 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 10214 17978
rect 10266 17926 10278 17978
rect 10330 17926 10342 17978
rect 10394 17926 10406 17978
rect 10458 17926 10470 17978
rect 10522 17926 16214 17978
rect 16266 17926 16278 17978
rect 16330 17926 16342 17978
rect 16394 17926 16406 17978
rect 16458 17926 16470 17978
rect 16522 17926 20792 17978
rect 1104 17904 20792 17926
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 13446 17864 13452 17876
rect 12676 17836 13452 17864
rect 12676 17824 12682 17836
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 14737 17867 14795 17873
rect 14737 17833 14749 17867
rect 14783 17864 14795 17867
rect 15470 17864 15476 17876
rect 14783 17836 15476 17864
rect 14783 17833 14795 17836
rect 14737 17827 14795 17833
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 18046 17824 18052 17876
rect 18104 17864 18110 17876
rect 19245 17867 19303 17873
rect 19245 17864 19257 17867
rect 18104 17836 19257 17864
rect 18104 17824 18110 17836
rect 19245 17833 19257 17836
rect 19291 17833 19303 17867
rect 19245 17827 19303 17833
rect 19610 17824 19616 17876
rect 19668 17824 19674 17876
rect 17773 17799 17831 17805
rect 17773 17765 17785 17799
rect 17819 17796 17831 17799
rect 18598 17796 18604 17808
rect 17819 17768 18604 17796
rect 17819 17765 17831 17768
rect 17773 17759 17831 17765
rect 18598 17756 18604 17768
rect 18656 17756 18662 17808
rect 5261 17731 5319 17737
rect 5261 17697 5273 17731
rect 5307 17728 5319 17731
rect 6086 17728 6092 17740
rect 5307 17700 6092 17728
rect 5307 17697 5319 17700
rect 5261 17691 5319 17697
rect 1670 17620 1676 17672
rect 1728 17660 1734 17672
rect 3237 17663 3295 17669
rect 3237 17660 3249 17663
rect 1728 17632 3249 17660
rect 1728 17620 1734 17632
rect 3237 17629 3249 17632
rect 3283 17660 3295 17663
rect 3283 17632 3648 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 2682 17552 2688 17604
rect 2740 17592 2746 17604
rect 2970 17595 3028 17601
rect 2970 17592 2982 17595
rect 2740 17564 2982 17592
rect 2740 17552 2746 17564
rect 2970 17561 2982 17564
rect 3016 17561 3028 17595
rect 2970 17555 3028 17561
rect 1394 17484 1400 17536
rect 1452 17524 1458 17536
rect 3620 17533 3648 17632
rect 3786 17620 3792 17672
rect 3844 17620 3850 17672
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 4479 17632 4537 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4525 17629 4537 17632
rect 4571 17629 4583 17663
rect 4525 17623 4583 17629
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17629 4767 17663
rect 4709 17623 4767 17629
rect 4724 17592 4752 17623
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 4893 17663 4951 17669
rect 4893 17660 4905 17663
rect 4856 17632 4905 17660
rect 4856 17620 4862 17632
rect 4893 17629 4905 17632
rect 4939 17629 4951 17663
rect 4893 17623 4951 17629
rect 5077 17663 5135 17669
rect 5077 17629 5089 17663
rect 5123 17629 5135 17663
rect 5077 17623 5135 17629
rect 5092 17592 5120 17623
rect 5350 17620 5356 17672
rect 5408 17620 5414 17672
rect 5552 17669 5580 17700
rect 6086 17688 6092 17700
rect 6144 17688 6150 17740
rect 16114 17688 16120 17740
rect 16172 17688 16178 17740
rect 17865 17731 17923 17737
rect 17865 17697 17877 17731
rect 17911 17728 17923 17731
rect 17954 17728 17960 17740
rect 17911 17700 17960 17728
rect 17911 17697 17923 17700
rect 17865 17691 17923 17697
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17728 19671 17731
rect 19978 17728 19984 17740
rect 19659 17700 19984 17728
rect 19659 17697 19671 17700
rect 19613 17691 19671 17697
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 5537 17663 5595 17669
rect 5537 17629 5549 17663
rect 5583 17629 5595 17663
rect 5537 17623 5595 17629
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 11514 17660 11520 17672
rect 9999 17632 11520 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 11514 17620 11520 17632
rect 11572 17660 11578 17672
rect 12989 17663 13047 17669
rect 12989 17660 13001 17663
rect 11572 17632 13001 17660
rect 11572 17620 11578 17632
rect 12989 17629 13001 17632
rect 13035 17660 13047 17663
rect 13722 17660 13728 17672
rect 13035 17632 13728 17660
rect 13035 17629 13047 17632
rect 12989 17623 13047 17629
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 15838 17620 15844 17672
rect 15896 17669 15902 17672
rect 15896 17660 15908 17669
rect 15896 17632 15941 17660
rect 15896 17623 15908 17632
rect 15896 17620 15902 17623
rect 16942 17620 16948 17672
rect 17000 17660 17006 17672
rect 17589 17663 17647 17669
rect 17589 17660 17601 17663
rect 17000 17632 17601 17660
rect 17000 17620 17006 17632
rect 17589 17629 17601 17632
rect 17635 17629 17647 17663
rect 17589 17623 17647 17629
rect 19426 17620 19432 17672
rect 19484 17620 19490 17672
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17660 19763 17663
rect 19794 17660 19800 17672
rect 19751 17632 19800 17660
rect 19751 17629 19763 17632
rect 19705 17623 19763 17629
rect 19794 17620 19800 17632
rect 19852 17620 19858 17672
rect 4724 17564 5120 17592
rect 5092 17536 5120 17564
rect 10220 17595 10278 17601
rect 10220 17561 10232 17595
rect 10266 17592 10278 17595
rect 10266 17564 11652 17592
rect 10266 17561 10278 17564
rect 10220 17555 10278 17561
rect 11624 17536 11652 17564
rect 12526 17552 12532 17604
rect 12584 17592 12590 17604
rect 12722 17595 12780 17601
rect 12722 17592 12734 17595
rect 12584 17564 12734 17592
rect 12584 17552 12590 17564
rect 12722 17561 12734 17564
rect 12768 17561 12780 17595
rect 12722 17555 12780 17561
rect 12894 17552 12900 17604
rect 12952 17592 12958 17604
rect 13081 17595 13139 17601
rect 13081 17592 13093 17595
rect 12952 17564 13093 17592
rect 12952 17552 12958 17564
rect 13081 17561 13093 17564
rect 13127 17561 13139 17595
rect 13081 17555 13139 17561
rect 13170 17552 13176 17604
rect 13228 17592 13234 17604
rect 13357 17595 13415 17601
rect 13357 17592 13369 17595
rect 13228 17564 13369 17592
rect 13228 17552 13234 17564
rect 13357 17561 13369 17564
rect 13403 17561 13415 17595
rect 13357 17555 13415 17561
rect 13446 17552 13452 17604
rect 13504 17552 13510 17604
rect 14274 17552 14280 17604
rect 14332 17592 14338 17604
rect 17957 17595 18015 17601
rect 17957 17592 17969 17595
rect 14332 17564 17969 17592
rect 14332 17552 14338 17564
rect 17957 17561 17969 17564
rect 18003 17592 18015 17595
rect 18046 17592 18052 17604
rect 18003 17564 18052 17592
rect 18003 17561 18015 17564
rect 17957 17555 18015 17561
rect 18046 17552 18052 17564
rect 18104 17552 18110 17604
rect 1857 17527 1915 17533
rect 1857 17524 1869 17527
rect 1452 17496 1869 17524
rect 1452 17484 1458 17496
rect 1857 17493 1869 17496
rect 1903 17493 1915 17527
rect 1857 17487 1915 17493
rect 3605 17527 3663 17533
rect 3605 17493 3617 17527
rect 3651 17524 3663 17527
rect 4246 17524 4252 17536
rect 3651 17496 4252 17524
rect 3651 17493 3663 17496
rect 3605 17487 3663 17493
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 4614 17484 4620 17536
rect 4672 17484 4678 17536
rect 5074 17484 5080 17536
rect 5132 17484 5138 17536
rect 5445 17527 5503 17533
rect 5445 17493 5457 17527
rect 5491 17524 5503 17527
rect 5534 17524 5540 17536
rect 5491 17496 5540 17524
rect 5491 17493 5503 17496
rect 5445 17487 5503 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 5626 17484 5632 17536
rect 5684 17484 5690 17536
rect 11333 17527 11391 17533
rect 11333 17493 11345 17527
rect 11379 17524 11391 17527
rect 11422 17524 11428 17536
rect 11379 17496 11428 17524
rect 11379 17493 11391 17496
rect 11333 17487 11391 17493
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 11606 17484 11612 17536
rect 11664 17484 11670 17536
rect 12986 17484 12992 17536
rect 13044 17524 13050 17536
rect 13265 17527 13323 17533
rect 13265 17524 13277 17527
rect 13044 17496 13277 17524
rect 13044 17484 13050 17496
rect 13265 17493 13277 17496
rect 13311 17493 13323 17527
rect 13265 17487 13323 17493
rect 13538 17484 13544 17536
rect 13596 17524 13602 17536
rect 13633 17527 13691 17533
rect 13633 17524 13645 17527
rect 13596 17496 13645 17524
rect 13596 17484 13602 17496
rect 13633 17493 13645 17496
rect 13679 17493 13691 17527
rect 13633 17487 13691 17493
rect 17678 17484 17684 17536
rect 17736 17484 17742 17536
rect 1104 17434 20792 17456
rect 1104 17382 7214 17434
rect 7266 17382 7278 17434
rect 7330 17382 7342 17434
rect 7394 17382 7406 17434
rect 7458 17382 7470 17434
rect 7522 17382 13214 17434
rect 13266 17382 13278 17434
rect 13330 17382 13342 17434
rect 13394 17382 13406 17434
rect 13458 17382 13470 17434
rect 13522 17382 19214 17434
rect 19266 17382 19278 17434
rect 19330 17382 19342 17434
rect 19394 17382 19406 17434
rect 19458 17382 19470 17434
rect 19522 17382 20792 17434
rect 1104 17360 20792 17382
rect 1670 17280 1676 17332
rect 1728 17280 1734 17332
rect 2682 17280 2688 17332
rect 2740 17280 2746 17332
rect 4614 17280 4620 17332
rect 4672 17280 4678 17332
rect 6656 17292 6960 17320
rect 4004 17255 4062 17261
rect 4004 17221 4016 17255
rect 4050 17252 4062 17255
rect 4632 17252 4660 17280
rect 4050 17224 4660 17252
rect 4050 17221 4062 17224
rect 4004 17215 4062 17221
rect 6656 17196 6684 17292
rect 6932 17252 6960 17292
rect 12894 17280 12900 17332
rect 12952 17280 12958 17332
rect 12986 17280 12992 17332
rect 13044 17280 13050 17332
rect 17037 17323 17095 17329
rect 17037 17289 17049 17323
rect 17083 17320 17095 17323
rect 17083 17292 18000 17320
rect 17083 17289 17095 17292
rect 17037 17283 17095 17289
rect 6932 17224 7590 17252
rect 11422 17212 11428 17264
rect 11480 17252 11486 17264
rect 12912 17252 12940 17280
rect 11480 17224 12940 17252
rect 11480 17212 11486 17224
rect 1394 17144 1400 17196
rect 1452 17184 1458 17196
rect 1765 17187 1823 17193
rect 1765 17184 1777 17187
rect 1452 17156 1777 17184
rect 1452 17144 1458 17156
rect 1765 17153 1777 17156
rect 1811 17153 1823 17187
rect 1765 17147 1823 17153
rect 5626 17144 5632 17196
rect 5684 17144 5690 17196
rect 5718 17144 5724 17196
rect 5776 17184 5782 17196
rect 6638 17184 6644 17196
rect 5776 17156 6644 17184
rect 5776 17144 5782 17156
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 6822 17144 6828 17196
rect 6880 17144 6886 17196
rect 9309 17187 9367 17193
rect 9309 17153 9321 17187
rect 9355 17184 9367 17187
rect 10229 17187 10287 17193
rect 10229 17184 10241 17187
rect 9355 17156 10241 17184
rect 9355 17153 9367 17156
rect 9309 17147 9367 17153
rect 10229 17153 10241 17156
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 11606 17144 11612 17196
rect 11664 17184 11670 17196
rect 11664 17156 12434 17184
rect 11664 17144 11670 17156
rect 1857 17119 1915 17125
rect 1857 17085 1869 17119
rect 1903 17116 1915 17119
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1903 17088 2053 17116
rect 1903 17085 1915 17088
rect 1857 17079 1915 17085
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 4246 17076 4252 17128
rect 4304 17076 4310 17128
rect 4338 17076 4344 17128
rect 4396 17076 4402 17128
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17116 4675 17119
rect 5644 17116 5672 17144
rect 4663 17088 5672 17116
rect 7101 17119 7159 17125
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 7101 17085 7113 17119
rect 7147 17116 7159 17119
rect 7650 17116 7656 17128
rect 7147 17088 7656 17116
rect 7147 17085 7159 17088
rect 7101 17079 7159 17085
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17116 9459 17119
rect 10134 17116 10140 17128
rect 9447 17088 10140 17116
rect 9447 17085 9459 17088
rect 9401 17079 9459 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 2869 16983 2927 16989
rect 2869 16949 2881 16983
rect 2915 16980 2927 16983
rect 3510 16980 3516 16992
rect 2915 16952 3516 16980
rect 2915 16949 2927 16952
rect 2869 16943 2927 16949
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 4264 16980 4292 17076
rect 5258 16980 5264 16992
rect 4264 16952 5264 16980
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 6089 16983 6147 16989
rect 6089 16949 6101 16983
rect 6135 16980 6147 16983
rect 6178 16980 6184 16992
rect 6135 16952 6184 16980
rect 6135 16949 6147 16952
rect 6089 16943 6147 16949
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 8570 16940 8576 16992
rect 8628 16940 8634 16992
rect 9582 16940 9588 16992
rect 9640 16940 9646 16992
rect 12406 16980 12434 17156
rect 12526 17144 12532 17196
rect 12584 17144 12590 17196
rect 12618 17144 12624 17196
rect 12676 17144 12682 17196
rect 12912 17193 12940 17224
rect 12897 17187 12955 17193
rect 12897 17153 12909 17187
rect 12943 17153 12955 17187
rect 12897 17147 12955 17153
rect 12544 17116 12572 17144
rect 12713 17119 12771 17125
rect 12713 17116 12725 17119
rect 12544 17088 12725 17116
rect 12713 17085 12725 17088
rect 12759 17085 12771 17119
rect 12713 17079 12771 17085
rect 12897 16983 12955 16989
rect 12897 16980 12909 16983
rect 12406 16952 12909 16980
rect 12897 16949 12909 16952
rect 12943 16980 12955 16983
rect 13004 16980 13032 17280
rect 17972 17264 18000 17292
rect 13078 17212 13084 17264
rect 13136 17252 13142 17264
rect 13265 17255 13323 17261
rect 13265 17252 13277 17255
rect 13136 17224 13277 17252
rect 13136 17212 13142 17224
rect 13265 17221 13277 17224
rect 13311 17221 13323 17255
rect 13265 17215 13323 17221
rect 13481 17255 13539 17261
rect 13481 17221 13493 17255
rect 13527 17252 13539 17255
rect 13630 17252 13636 17264
rect 13527 17224 13636 17252
rect 13527 17221 13539 17224
rect 13481 17215 13539 17221
rect 13630 17212 13636 17224
rect 13688 17212 13694 17264
rect 17954 17212 17960 17264
rect 18012 17212 18018 17264
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17184 13783 17187
rect 13906 17184 13912 17196
rect 13771 17156 13912 17184
rect 13771 17153 13783 17156
rect 13725 17147 13783 17153
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 14458 17144 14464 17196
rect 14516 17144 14522 17196
rect 18161 17187 18219 17193
rect 18161 17153 18173 17187
rect 18207 17184 18219 17187
rect 18690 17184 18696 17196
rect 18207 17156 18696 17184
rect 18207 17153 18219 17156
rect 18161 17147 18219 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 19236 17187 19294 17193
rect 19236 17153 19248 17187
rect 19282 17184 19294 17187
rect 19610 17184 19616 17196
rect 19282 17156 19616 17184
rect 19282 17153 19294 17156
rect 19236 17147 19294 17153
rect 19610 17144 19616 17156
rect 19668 17144 19674 17196
rect 13817 17119 13875 17125
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 14476 17116 14504 17144
rect 13863 17088 14504 17116
rect 18417 17119 18475 17125
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 18417 17085 18429 17119
rect 18463 17116 18475 17119
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 18463 17088 18981 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 18969 17085 18981 17088
rect 19015 17085 19027 17119
rect 18969 17079 19027 17085
rect 13081 17051 13139 17057
rect 13081 17017 13093 17051
rect 13127 17048 13139 17051
rect 13127 17020 13860 17048
rect 13127 17017 13139 17020
rect 13081 17011 13139 17017
rect 12943 16952 13032 16980
rect 13449 16983 13507 16989
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 13449 16949 13461 16983
rect 13495 16980 13507 16983
rect 13538 16980 13544 16992
rect 13495 16952 13544 16980
rect 13495 16949 13507 16952
rect 13449 16943 13507 16949
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 13633 16983 13691 16989
rect 13633 16949 13645 16983
rect 13679 16980 13691 16983
rect 13722 16980 13728 16992
rect 13679 16952 13728 16980
rect 13679 16949 13691 16952
rect 13633 16943 13691 16949
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 13832 16989 13860 17020
rect 13817 16983 13875 16989
rect 13817 16949 13829 16983
rect 13863 16949 13875 16983
rect 13817 16943 13875 16949
rect 14090 16940 14096 16992
rect 14148 16940 14154 16992
rect 18138 16940 18144 16992
rect 18196 16980 18202 16992
rect 18432 16980 18460 17079
rect 18196 16952 18460 16980
rect 20349 16983 20407 16989
rect 18196 16940 18202 16952
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20395 16952 20852 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 1104 16890 20792 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 10214 16890
rect 10266 16838 10278 16890
rect 10330 16838 10342 16890
rect 10394 16838 10406 16890
rect 10458 16838 10470 16890
rect 10522 16838 16214 16890
rect 16266 16838 16278 16890
rect 16330 16838 16342 16890
rect 16394 16838 16406 16890
rect 16458 16838 16470 16890
rect 16522 16838 20792 16890
rect 1104 16816 20792 16838
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 6178 16785 6184 16788
rect 3973 16779 4031 16785
rect 3973 16776 3985 16779
rect 3936 16748 3985 16776
rect 3936 16736 3942 16748
rect 3973 16745 3985 16748
rect 4019 16745 4031 16779
rect 3973 16739 4031 16745
rect 6168 16779 6184 16785
rect 6168 16745 6180 16779
rect 6168 16739 6184 16745
rect 6178 16736 6184 16739
rect 6236 16736 6242 16788
rect 7650 16736 7656 16788
rect 7708 16736 7714 16788
rect 10134 16776 10140 16788
rect 8588 16748 10140 16776
rect 8588 16708 8616 16748
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10594 16736 10600 16788
rect 10652 16776 10658 16788
rect 10870 16776 10876 16788
rect 10652 16748 10876 16776
rect 10652 16736 10658 16748
rect 10870 16736 10876 16748
rect 10928 16776 10934 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 10928 16748 11069 16776
rect 10928 16736 10934 16748
rect 11057 16745 11069 16748
rect 11103 16745 11115 16779
rect 11057 16739 11115 16745
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 13780 16748 15792 16776
rect 13780 16736 13786 16748
rect 8496 16680 8616 16708
rect 14921 16711 14979 16717
rect 1673 16643 1731 16649
rect 1673 16609 1685 16643
rect 1719 16640 1731 16643
rect 2038 16640 2044 16652
rect 1719 16612 2044 16640
rect 1719 16609 1731 16612
rect 1673 16603 1731 16609
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 5813 16643 5871 16649
rect 5813 16609 5825 16643
rect 5859 16640 5871 16643
rect 5859 16612 7420 16640
rect 5859 16609 5871 16612
rect 5813 16603 5871 16609
rect 3329 16575 3387 16581
rect 3329 16541 3341 16575
rect 3375 16572 3387 16575
rect 5258 16572 5264 16584
rect 3375 16544 5264 16572
rect 3375 16541 3387 16544
rect 3329 16535 3387 16541
rect 5258 16532 5264 16544
rect 5316 16572 5322 16584
rect 5828 16572 5856 16603
rect 5316 16544 5856 16572
rect 5905 16575 5963 16581
rect 5316 16532 5322 16544
rect 5905 16541 5917 16575
rect 5951 16541 5963 16575
rect 7392 16572 7420 16612
rect 8496 16581 8524 16680
rect 14921 16677 14933 16711
rect 14967 16708 14979 16711
rect 14967 16680 15700 16708
rect 14967 16677 14979 16680
rect 14921 16671 14979 16677
rect 9306 16640 9312 16652
rect 8680 16612 9312 16640
rect 8680 16584 8708 16612
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 14274 16600 14280 16652
rect 14332 16640 14338 16652
rect 14332 16612 15056 16640
rect 14332 16600 14338 16612
rect 8481 16575 8539 16581
rect 7392 16544 8248 16572
rect 5905 16535 5963 16541
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 1489 16507 1547 16513
rect 1489 16504 1501 16507
rect 992 16476 1501 16504
rect 992 16464 998 16476
rect 1489 16473 1501 16476
rect 1535 16473 1547 16507
rect 1489 16467 1547 16473
rect 2682 16464 2688 16516
rect 2740 16504 2746 16516
rect 3062 16507 3120 16513
rect 3062 16504 3074 16507
rect 2740 16476 3074 16504
rect 2740 16464 2746 16476
rect 3062 16473 3074 16476
rect 3108 16473 3120 16507
rect 3789 16507 3847 16513
rect 3789 16504 3801 16507
rect 3062 16467 3120 16473
rect 3436 16476 3801 16504
rect 3436 16448 3464 16476
rect 3789 16473 3801 16476
rect 3835 16473 3847 16507
rect 5074 16504 5080 16516
rect 3789 16467 3847 16473
rect 4172 16476 5080 16504
rect 1670 16396 1676 16448
rect 1728 16436 1734 16448
rect 1949 16439 2007 16445
rect 1949 16436 1961 16439
rect 1728 16408 1961 16436
rect 1728 16396 1734 16408
rect 1949 16405 1961 16408
rect 1995 16436 2007 16439
rect 3326 16436 3332 16448
rect 1995 16408 3332 16436
rect 1995 16405 2007 16408
rect 1949 16399 2007 16405
rect 3326 16396 3332 16408
rect 3384 16396 3390 16448
rect 3418 16396 3424 16448
rect 3476 16396 3482 16448
rect 3510 16396 3516 16448
rect 3568 16436 3574 16448
rect 4172 16445 4200 16476
rect 5074 16464 5080 16476
rect 5132 16464 5138 16516
rect 5534 16464 5540 16516
rect 5592 16513 5598 16516
rect 5592 16504 5604 16513
rect 5592 16476 5637 16504
rect 5592 16467 5604 16476
rect 5592 16464 5598 16467
rect 3989 16439 4047 16445
rect 3989 16436 4001 16439
rect 3568 16408 4001 16436
rect 3568 16396 3574 16408
rect 3989 16405 4001 16408
rect 4035 16405 4047 16439
rect 3989 16399 4047 16405
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16405 4215 16439
rect 4157 16399 4215 16405
rect 4433 16439 4491 16445
rect 4433 16405 4445 16439
rect 4479 16436 4491 16439
rect 4614 16436 4620 16448
rect 4479 16408 4620 16436
rect 4479 16405 4491 16408
rect 4433 16399 4491 16405
rect 4614 16396 4620 16408
rect 4672 16436 4678 16448
rect 4890 16436 4896 16448
rect 4672 16408 4896 16436
rect 4672 16396 4678 16408
rect 4890 16396 4896 16408
rect 4948 16436 4954 16448
rect 5920 16436 5948 16535
rect 6638 16464 6644 16516
rect 6696 16464 6702 16516
rect 6822 16436 6828 16448
rect 4948 16408 6828 16436
rect 4948 16396 4954 16408
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 8220 16445 8248 16544
rect 8481 16541 8493 16575
rect 8527 16541 8539 16575
rect 8481 16535 8539 16541
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16541 8631 16575
rect 8573 16535 8631 16541
rect 8588 16504 8616 16535
rect 8662 16532 8668 16584
rect 8720 16532 8726 16584
rect 8757 16575 8815 16581
rect 8757 16541 8769 16575
rect 8803 16572 8815 16575
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 8803 16544 9137 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 9125 16541 9137 16544
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 11146 16532 11152 16584
rect 11204 16532 11210 16584
rect 11422 16581 11428 16584
rect 11416 16572 11428 16581
rect 11383 16544 11428 16572
rect 11416 16535 11428 16544
rect 11422 16532 11428 16535
rect 11480 16532 11486 16584
rect 14090 16532 14096 16584
rect 14148 16572 14154 16584
rect 14921 16575 14979 16581
rect 14921 16572 14933 16575
rect 14148 16544 14933 16572
rect 14148 16532 14154 16544
rect 14921 16541 14933 16544
rect 14967 16541 14979 16575
rect 15028 16572 15056 16612
rect 15102 16600 15108 16652
rect 15160 16600 15166 16652
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16640 15255 16643
rect 15470 16640 15476 16652
rect 15243 16612 15476 16640
rect 15243 16609 15255 16612
rect 15197 16603 15255 16609
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15562 16600 15568 16652
rect 15620 16600 15626 16652
rect 15289 16575 15347 16581
rect 15289 16572 15301 16575
rect 15028 16544 15301 16572
rect 14921 16535 14979 16541
rect 15289 16541 15301 16544
rect 15335 16572 15347 16575
rect 15381 16575 15439 16581
rect 15381 16572 15393 16575
rect 15335 16544 15393 16572
rect 15335 16541 15347 16544
rect 15289 16535 15347 16541
rect 15381 16541 15393 16544
rect 15427 16541 15439 16575
rect 15672 16572 15700 16680
rect 15764 16649 15792 16748
rect 18598 16736 18604 16788
rect 18656 16736 18662 16788
rect 18690 16736 18696 16788
rect 18748 16736 18754 16788
rect 19061 16779 19119 16785
rect 19061 16745 19073 16779
rect 19107 16776 19119 16779
rect 19610 16776 19616 16788
rect 19107 16748 19616 16776
rect 19107 16745 19119 16748
rect 19061 16739 19119 16745
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 16025 16643 16083 16649
rect 16025 16609 16037 16643
rect 16071 16640 16083 16643
rect 17310 16640 17316 16652
rect 16071 16612 17316 16640
rect 16071 16609 16083 16612
rect 16025 16603 16083 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 17586 16600 17592 16652
rect 17644 16640 17650 16652
rect 17865 16643 17923 16649
rect 17865 16640 17877 16643
rect 17644 16612 17877 16640
rect 17644 16600 17650 16612
rect 17865 16609 17877 16612
rect 17911 16609 17923 16643
rect 17865 16603 17923 16609
rect 18049 16643 18107 16649
rect 18049 16609 18061 16643
rect 18095 16640 18107 16643
rect 18708 16640 18736 16736
rect 19797 16711 19855 16717
rect 19797 16677 19809 16711
rect 19843 16708 19855 16711
rect 20824 16708 20852 16952
rect 19843 16680 20852 16708
rect 19843 16677 19855 16680
rect 19797 16671 19855 16677
rect 19812 16640 19840 16671
rect 18095 16612 18644 16640
rect 18708 16612 19840 16640
rect 18095 16609 18107 16612
rect 18049 16603 18107 16609
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15672 16544 15853 16572
rect 15381 16535 15439 16541
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 17773 16575 17831 16581
rect 17773 16572 17785 16575
rect 17736 16544 17785 16572
rect 17736 16532 17742 16544
rect 17773 16541 17785 16544
rect 17819 16541 17831 16575
rect 17773 16535 17831 16541
rect 17954 16532 17960 16584
rect 18012 16572 18018 16584
rect 18141 16575 18199 16581
rect 18141 16572 18153 16575
rect 18012 16544 18153 16572
rect 18012 16532 18018 16544
rect 18141 16541 18153 16544
rect 18187 16541 18199 16575
rect 18141 16535 18199 16541
rect 9674 16504 9680 16516
rect 8588 16476 9680 16504
rect 9674 16464 9680 16476
rect 9732 16464 9738 16516
rect 11882 16504 11888 16516
rect 10810 16476 11888 16504
rect 11882 16464 11888 16476
rect 11940 16504 11946 16516
rect 11940 16476 14228 16504
rect 11940 16464 11946 16476
rect 8205 16439 8263 16445
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 8294 16436 8300 16448
rect 8251 16408 8300 16436
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 8294 16396 8300 16408
rect 8352 16436 8358 16448
rect 8662 16436 8668 16448
rect 8352 16408 8668 16436
rect 8352 16396 8358 16408
rect 8662 16396 8668 16408
rect 8720 16396 8726 16448
rect 8938 16396 8944 16448
rect 8996 16396 9002 16448
rect 12526 16396 12532 16448
rect 12584 16396 12590 16448
rect 14200 16436 14228 16476
rect 17586 16464 17592 16516
rect 17644 16464 17650 16516
rect 18046 16464 18052 16516
rect 18104 16504 18110 16516
rect 18233 16507 18291 16513
rect 18233 16504 18245 16507
rect 18104 16476 18245 16504
rect 18104 16464 18110 16476
rect 18233 16473 18245 16476
rect 18279 16473 18291 16507
rect 18233 16467 18291 16473
rect 14918 16436 14924 16448
rect 14200 16408 14924 16436
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 18616 16436 18644 16612
rect 18800 16581 18828 16612
rect 18785 16575 18843 16581
rect 18785 16541 18797 16575
rect 18831 16541 18843 16575
rect 18785 16535 18843 16541
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19521 16575 19579 16581
rect 19521 16572 19533 16575
rect 18923 16544 19533 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 18984 16516 19012 16544
rect 19521 16541 19533 16544
rect 19567 16541 19579 16575
rect 19702 16572 19708 16584
rect 19521 16535 19579 16541
rect 19628 16544 19708 16572
rect 18966 16464 18972 16516
rect 19024 16464 19030 16516
rect 19058 16464 19064 16516
rect 19116 16504 19122 16516
rect 19429 16507 19487 16513
rect 19429 16504 19441 16507
rect 19116 16476 19441 16504
rect 19116 16464 19122 16476
rect 19429 16473 19441 16476
rect 19475 16504 19487 16507
rect 19628 16504 19656 16544
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 19475 16476 19656 16504
rect 19475 16473 19487 16476
rect 19429 16467 19487 16473
rect 19245 16439 19303 16445
rect 19245 16436 19257 16439
rect 18616 16408 19257 16436
rect 19245 16405 19257 16408
rect 19291 16405 19303 16439
rect 19245 16399 19303 16405
rect 19610 16396 19616 16448
rect 19668 16396 19674 16448
rect 1104 16346 20792 16368
rect 1104 16294 7214 16346
rect 7266 16294 7278 16346
rect 7330 16294 7342 16346
rect 7394 16294 7406 16346
rect 7458 16294 7470 16346
rect 7522 16294 13214 16346
rect 13266 16294 13278 16346
rect 13330 16294 13342 16346
rect 13394 16294 13406 16346
rect 13458 16294 13470 16346
rect 13522 16294 19214 16346
rect 19266 16294 19278 16346
rect 19330 16294 19342 16346
rect 19394 16294 19406 16346
rect 19458 16294 19470 16346
rect 19522 16294 20792 16346
rect 1104 16272 20792 16294
rect 2682 16192 2688 16244
rect 2740 16192 2746 16244
rect 3237 16235 3295 16241
rect 3237 16201 3249 16235
rect 3283 16232 3295 16235
rect 4249 16235 4307 16241
rect 4249 16232 4261 16235
rect 3283 16204 4261 16232
rect 3283 16201 3295 16204
rect 3237 16195 3295 16201
rect 4249 16201 4261 16204
rect 4295 16232 4307 16235
rect 5258 16232 5264 16244
rect 4295 16204 5264 16232
rect 4295 16201 4307 16204
rect 4249 16195 4307 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 5350 16192 5356 16244
rect 5408 16192 5414 16244
rect 8938 16232 8944 16244
rect 8128 16204 8944 16232
rect 3418 16164 3424 16176
rect 2746 16136 3424 16164
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 1452 16068 1593 16096
rect 1452 16056 1458 16068
rect 1581 16065 1593 16068
rect 1627 16096 1639 16099
rect 2746 16096 2774 16136
rect 3418 16124 3424 16136
rect 3476 16124 3482 16176
rect 3510 16124 3516 16176
rect 3568 16164 3574 16176
rect 3605 16167 3663 16173
rect 3605 16164 3617 16167
rect 3568 16136 3617 16164
rect 3568 16124 3574 16136
rect 3605 16133 3617 16136
rect 3651 16133 3663 16167
rect 3605 16127 3663 16133
rect 4985 16167 5043 16173
rect 4985 16133 4997 16167
rect 5031 16164 5043 16167
rect 5368 16164 5396 16192
rect 8128 16173 8156 16204
rect 8938 16192 8944 16204
rect 8996 16192 9002 16244
rect 9585 16235 9643 16241
rect 9585 16201 9597 16235
rect 9631 16201 9643 16235
rect 9585 16195 9643 16201
rect 5031 16136 5396 16164
rect 8113 16167 8171 16173
rect 5031 16133 5043 16136
rect 4985 16127 5043 16133
rect 8113 16133 8125 16167
rect 8159 16133 8171 16167
rect 8113 16127 8171 16133
rect 8846 16124 8852 16176
rect 8904 16124 8910 16176
rect 9600 16164 9628 16195
rect 9674 16192 9680 16244
rect 9732 16192 9738 16244
rect 10134 16192 10140 16244
rect 10192 16192 10198 16244
rect 14921 16235 14979 16241
rect 14921 16201 14933 16235
rect 14967 16232 14979 16235
rect 15102 16232 15108 16244
rect 14967 16204 15108 16232
rect 14967 16201 14979 16204
rect 14921 16195 14979 16201
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 15528 16204 16773 16232
rect 15528 16192 15534 16204
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 16761 16195 16819 16201
rect 19610 16192 19616 16244
rect 19668 16232 19674 16244
rect 19981 16235 20039 16241
rect 19981 16232 19993 16235
rect 19668 16204 19993 16232
rect 19668 16192 19674 16204
rect 19981 16201 19993 16204
rect 20027 16201 20039 16235
rect 19981 16195 20039 16201
rect 9861 16167 9919 16173
rect 9861 16164 9873 16167
rect 9600 16136 9873 16164
rect 9861 16133 9873 16136
rect 9907 16164 9919 16167
rect 18868 16167 18926 16173
rect 9907 16136 10180 16164
rect 9907 16133 9919 16136
rect 9861 16127 9919 16133
rect 10152 16108 10180 16136
rect 14752 16136 16436 16164
rect 1627 16068 2774 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 3326 16056 3332 16108
rect 3384 16056 3390 16108
rect 4890 16056 4896 16108
rect 4948 16056 4954 16108
rect 5074 16056 5080 16108
rect 5132 16056 5138 16108
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 10045 16099 10103 16105
rect 10045 16096 10057 16099
rect 9824 16068 10057 16096
rect 9824 16056 9830 16068
rect 10045 16065 10057 16068
rect 10091 16065 10103 16099
rect 10045 16059 10103 16065
rect 1670 15988 1676 16040
rect 1728 15988 1734 16040
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1995 16000 2053 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 3344 16028 3372 16056
rect 3878 16028 3884 16040
rect 3344 16000 3884 16028
rect 2041 15991 2099 15997
rect 3878 15988 3884 16000
rect 3936 15988 3942 16040
rect 7837 16031 7895 16037
rect 7837 15997 7849 16031
rect 7883 15997 7895 16031
rect 10060 16028 10088 16059
rect 10134 16056 10140 16108
rect 10192 16056 10198 16108
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 10336 16028 10364 16059
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 14752 16105 14780 16136
rect 13153 16099 13211 16105
rect 13153 16096 13165 16099
rect 13044 16068 13165 16096
rect 13044 16056 13050 16068
rect 13153 16065 13165 16068
rect 13199 16065 13211 16099
rect 14461 16099 14519 16105
rect 14461 16096 14473 16099
rect 13153 16059 13211 16065
rect 14384 16068 14473 16096
rect 10060 16000 10364 16028
rect 7837 15991 7895 15997
rect 3605 15963 3663 15969
rect 3605 15929 3617 15963
rect 3651 15960 3663 15963
rect 3786 15960 3792 15972
rect 3651 15932 3792 15960
rect 3651 15929 3663 15932
rect 3605 15923 3663 15929
rect 3786 15920 3792 15932
rect 3844 15920 3850 15972
rect 7745 15895 7803 15901
rect 7745 15861 7757 15895
rect 7791 15892 7803 15895
rect 7852 15892 7880 15991
rect 12802 15988 12808 16040
rect 12860 16028 12866 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12860 16000 12909 16028
rect 12860 15988 12866 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 12897 15991 12955 15997
rect 14384 15904 14412 16068
rect 14461 16065 14473 16068
rect 14507 16065 14519 16099
rect 14461 16059 14519 16065
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 15269 16099 15327 16105
rect 15269 16096 15281 16099
rect 14737 16059 14795 16065
rect 14936 16068 15281 16096
rect 14642 15988 14648 16040
rect 14700 15988 14706 16040
rect 14936 16028 14964 16068
rect 15269 16065 15281 16068
rect 15315 16096 15327 16099
rect 15654 16096 15660 16108
rect 15315 16068 15660 16096
rect 15315 16065 15327 16068
rect 15269 16059 15327 16065
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 16408 16096 16436 16136
rect 18868 16133 18880 16167
rect 18914 16164 18926 16167
rect 18966 16164 18972 16176
rect 18914 16136 18972 16164
rect 18914 16133 18926 16136
rect 18868 16127 18926 16133
rect 18966 16124 18972 16136
rect 19024 16164 19030 16176
rect 19886 16164 19892 16176
rect 19024 16136 19892 16164
rect 19024 16124 19030 16136
rect 19886 16124 19892 16136
rect 19944 16124 19950 16176
rect 17874 16099 17932 16105
rect 17874 16096 17886 16099
rect 16408 16068 17886 16096
rect 14752 16000 14964 16028
rect 15013 16031 15071 16037
rect 7926 15892 7932 15904
rect 7791 15864 7932 15892
rect 7791 15861 7803 15864
rect 7745 15855 7803 15861
rect 7926 15852 7932 15864
rect 7984 15892 7990 15904
rect 8294 15892 8300 15904
rect 7984 15864 8300 15892
rect 7984 15852 7990 15864
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 14090 15892 14096 15904
rect 12492 15864 14096 15892
rect 12492 15852 12498 15864
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 14277 15895 14335 15901
rect 14277 15861 14289 15895
rect 14323 15892 14335 15895
rect 14366 15892 14372 15904
rect 14323 15864 14372 15892
rect 14323 15861 14335 15864
rect 14277 15855 14335 15861
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 14752 15901 14780 16000
rect 15013 15997 15025 16031
rect 15059 15997 15071 16031
rect 15013 15991 15071 15997
rect 14737 15895 14795 15901
rect 14737 15861 14749 15895
rect 14783 15861 14795 15895
rect 15028 15892 15056 15991
rect 16114 15920 16120 15972
rect 16172 15960 16178 15972
rect 16408 15969 16436 16068
rect 17874 16065 17886 16068
rect 17920 16065 17932 16099
rect 17874 16059 17932 16065
rect 18138 16056 18144 16108
rect 18196 16096 18202 16108
rect 18601 16099 18659 16105
rect 18601 16096 18613 16099
rect 18196 16068 18613 16096
rect 18196 16056 18202 16068
rect 18601 16065 18613 16068
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 16393 15963 16451 15969
rect 16393 15960 16405 15963
rect 16172 15932 16405 15960
rect 16172 15920 16178 15932
rect 16393 15929 16405 15932
rect 16439 15929 16451 15963
rect 16393 15923 16451 15929
rect 15286 15892 15292 15904
rect 15028 15864 15292 15892
rect 14737 15855 14795 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 17862 15892 17868 15904
rect 15436 15864 17868 15892
rect 15436 15852 15442 15864
rect 17862 15852 17868 15864
rect 17920 15852 17926 15904
rect 1104 15802 20792 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 10214 15802
rect 10266 15750 10278 15802
rect 10330 15750 10342 15802
rect 10394 15750 10406 15802
rect 10458 15750 10470 15802
rect 10522 15750 16214 15802
rect 16266 15750 16278 15802
rect 16330 15750 16342 15802
rect 16394 15750 16406 15802
rect 16458 15750 16470 15802
rect 16522 15750 20792 15802
rect 1104 15728 20792 15750
rect 12434 15688 12440 15700
rect 6840 15660 12440 15688
rect 3510 15580 3516 15632
rect 3568 15580 3574 15632
rect 6086 15580 6092 15632
rect 6144 15620 6150 15632
rect 6840 15629 6868 15660
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 12526 15648 12532 15700
rect 12584 15648 12590 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 12728 15660 13461 15688
rect 6825 15623 6883 15629
rect 6825 15620 6837 15623
rect 6144 15592 6837 15620
rect 6144 15580 6150 15592
rect 6825 15589 6837 15592
rect 6871 15589 6883 15623
rect 6825 15583 6883 15589
rect 1670 15444 1676 15496
rect 1728 15484 1734 15496
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1728 15456 2053 15484
rect 1728 15444 1734 15456
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 3528 15484 3556 15580
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 3528 15456 4169 15484
rect 2041 15447 2099 15453
rect 4157 15453 4169 15456
rect 4203 15453 4215 15487
rect 6932 15484 6960 15515
rect 11146 15512 11152 15564
rect 11204 15552 11210 15564
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 11204 15524 11253 15552
rect 11204 15512 11210 15524
rect 11241 15521 11253 15524
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 7193 15487 7251 15493
rect 7193 15484 7205 15487
rect 6932 15456 7205 15484
rect 4157 15447 4215 15453
rect 7193 15453 7205 15456
rect 7239 15453 7251 15487
rect 7193 15447 7251 15453
rect 6457 15419 6515 15425
rect 6457 15385 6469 15419
rect 6503 15416 6515 15419
rect 7834 15416 7840 15428
rect 6503 15388 7840 15416
rect 6503 15385 6515 15388
rect 6457 15379 6515 15385
rect 7834 15376 7840 15388
rect 7892 15376 7898 15428
rect 8846 15376 8852 15428
rect 8904 15416 8910 15428
rect 9858 15416 9864 15428
rect 8904 15388 9864 15416
rect 8904 15376 8910 15388
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 11508 15419 11566 15425
rect 11508 15385 11520 15419
rect 11554 15416 11566 15419
rect 12544 15416 12572 15648
rect 12728 15496 12756 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 13449 15651 13507 15657
rect 13630 15648 13636 15700
rect 13688 15648 13694 15700
rect 13906 15648 13912 15700
rect 13964 15648 13970 15700
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 14148 15660 15056 15688
rect 14148 15648 14154 15660
rect 12805 15623 12863 15629
rect 12805 15589 12817 15623
rect 12851 15620 12863 15623
rect 12986 15620 12992 15632
rect 12851 15592 12992 15620
rect 12851 15589 12863 15592
rect 12805 15583 12863 15589
rect 12986 15580 12992 15592
rect 13044 15580 13050 15632
rect 13357 15623 13415 15629
rect 13357 15589 13369 15623
rect 13403 15620 13415 15623
rect 13648 15620 13676 15648
rect 13403 15592 13676 15620
rect 15028 15620 15056 15660
rect 15562 15648 15568 15700
rect 15620 15688 15626 15700
rect 15657 15691 15715 15697
rect 15657 15688 15669 15691
rect 15620 15660 15669 15688
rect 15620 15648 15626 15660
rect 15657 15657 15669 15660
rect 15703 15657 15715 15691
rect 15657 15651 15715 15657
rect 16114 15648 16120 15700
rect 16172 15648 16178 15700
rect 16132 15620 16160 15648
rect 16209 15623 16267 15629
rect 16209 15620 16221 15623
rect 15028 15592 15608 15620
rect 16132 15592 16221 15620
rect 13403 15589 13415 15592
rect 13357 15583 13415 15589
rect 13004 15552 13032 15580
rect 15580 15552 15608 15592
rect 16209 15589 16221 15592
rect 16255 15589 16267 15623
rect 16209 15583 16267 15589
rect 18230 15580 18236 15632
rect 18288 15580 18294 15632
rect 18248 15552 18276 15580
rect 13004 15524 13768 15552
rect 15580 15524 18276 15552
rect 12710 15444 12716 15496
rect 12768 15484 12774 15496
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 12768 15456 13001 15484
rect 12768 15444 12774 15456
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 13078 15444 13084 15496
rect 13136 15484 13142 15496
rect 13740 15493 13768 15524
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 13136 15456 13645 15484
rect 13136 15444 13142 15456
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15484 14151 15487
rect 14182 15484 14188 15496
rect 14139 15456 14188 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 14366 15493 14372 15496
rect 14360 15447 14372 15493
rect 14424 15484 14430 15496
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 14424 15456 15853 15484
rect 14366 15444 14372 15447
rect 14424 15444 14430 15456
rect 15841 15453 15853 15456
rect 15887 15453 15899 15487
rect 15841 15447 15899 15453
rect 17310 15444 17316 15496
rect 17368 15444 17374 15496
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15484 17555 15487
rect 17586 15484 17592 15496
rect 17543 15456 17592 15484
rect 17543 15453 17555 15456
rect 17497 15447 17555 15453
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15484 17739 15487
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17727 15456 17785 15484
rect 17727 15453 17739 15456
rect 17681 15447 17739 15453
rect 17773 15453 17785 15456
rect 17819 15453 17831 15487
rect 17773 15447 17831 15453
rect 17862 15444 17868 15496
rect 17920 15484 17926 15496
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 17920 15456 18061 15484
rect 17920 15444 17926 15456
rect 18049 15453 18061 15456
rect 18095 15484 18107 15487
rect 20254 15484 20260 15496
rect 18095 15456 20260 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 13449 15419 13507 15425
rect 13449 15416 13461 15419
rect 11554 15388 13461 15416
rect 11554 15385 11566 15388
rect 11508 15379 11566 15385
rect 1854 15308 1860 15360
rect 1912 15348 1918 15360
rect 1949 15351 2007 15357
rect 1949 15348 1961 15351
rect 1912 15320 1961 15348
rect 1912 15308 1918 15320
rect 1949 15317 1961 15320
rect 1995 15317 2007 15351
rect 1949 15311 2007 15317
rect 4249 15351 4307 15357
rect 4249 15317 4261 15351
rect 4295 15348 4307 15351
rect 5994 15348 6000 15360
rect 4295 15320 6000 15348
rect 4295 15317 4307 15320
rect 4249 15311 4307 15317
rect 5994 15308 6000 15320
rect 6052 15308 6058 15360
rect 7006 15308 7012 15360
rect 7064 15308 7070 15360
rect 12526 15308 12532 15360
rect 12584 15348 12590 15360
rect 13188 15357 13216 15388
rect 13449 15385 13461 15388
rect 13495 15385 13507 15419
rect 13449 15379 13507 15385
rect 14642 15376 14648 15428
rect 14700 15376 14706 15428
rect 15933 15419 15991 15425
rect 15933 15416 15945 15419
rect 15488 15388 15945 15416
rect 12621 15351 12679 15357
rect 12621 15348 12633 15351
rect 12584 15320 12633 15348
rect 12584 15308 12590 15320
rect 12621 15317 12633 15320
rect 12667 15317 12679 15351
rect 12621 15311 12679 15317
rect 13173 15351 13231 15357
rect 13173 15317 13185 15351
rect 13219 15317 13231 15351
rect 14660 15348 14688 15376
rect 15488 15357 15516 15388
rect 15933 15385 15945 15388
rect 15979 15385 15991 15419
rect 15933 15379 15991 15385
rect 17129 15419 17187 15425
rect 17129 15385 17141 15419
rect 17175 15416 17187 15419
rect 17954 15416 17960 15428
rect 17175 15388 17960 15416
rect 17175 15385 17187 15388
rect 17129 15379 17187 15385
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 14660 15320 15485 15348
rect 13173 15311 13231 15317
rect 15473 15317 15485 15320
rect 15519 15317 15531 15351
rect 15473 15311 15531 15317
rect 15654 15308 15660 15360
rect 15712 15348 15718 15360
rect 16025 15351 16083 15357
rect 16025 15348 16037 15351
rect 15712 15320 16037 15348
rect 15712 15308 15718 15320
rect 16025 15317 16037 15320
rect 16071 15317 16083 15351
rect 16025 15311 16083 15317
rect 17405 15351 17463 15357
rect 17405 15317 17417 15351
rect 17451 15348 17463 15351
rect 18230 15348 18236 15360
rect 17451 15320 18236 15348
rect 17451 15317 17463 15320
rect 17405 15311 17463 15317
rect 18230 15308 18236 15320
rect 18288 15308 18294 15360
rect 1104 15258 20792 15280
rect 1104 15206 7214 15258
rect 7266 15206 7278 15258
rect 7330 15206 7342 15258
rect 7394 15206 7406 15258
rect 7458 15206 7470 15258
rect 7522 15206 13214 15258
rect 13266 15206 13278 15258
rect 13330 15206 13342 15258
rect 13394 15206 13406 15258
rect 13458 15206 13470 15258
rect 13522 15206 19214 15258
rect 19266 15206 19278 15258
rect 19330 15206 19342 15258
rect 19394 15206 19406 15258
rect 19458 15206 19470 15258
rect 19522 15206 20792 15258
rect 1104 15184 20792 15206
rect 1670 15104 1676 15156
rect 1728 15104 1734 15156
rect 7006 15144 7012 15156
rect 3436 15116 4108 15144
rect 1688 15076 1716 15104
rect 3436 15076 3464 15116
rect 1412 15048 1716 15076
rect 2898 15048 3464 15076
rect 1412 15017 1440 15048
rect 3510 15036 3516 15088
rect 3568 15076 3574 15088
rect 3786 15076 3792 15088
rect 3568 15048 3792 15076
rect 3568 15036 3574 15048
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 3878 15036 3884 15088
rect 3936 15036 3942 15088
rect 4080 15020 4108 15116
rect 6656 15116 7012 15144
rect 6656 15085 6684 15116
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 9824 15116 9873 15144
rect 9824 15104 9830 15116
rect 9861 15113 9873 15116
rect 9907 15113 9919 15147
rect 12710 15144 12716 15156
rect 9861 15107 9919 15113
rect 12360 15116 12716 15144
rect 6641 15079 6699 15085
rect 6641 15045 6653 15079
rect 6687 15045 6699 15079
rect 6641 15039 6699 15045
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 3326 14968 3332 15020
rect 3384 14968 3390 15020
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 1670 14900 1676 14952
rect 1728 14900 1734 14952
rect 3620 14940 3648 14971
rect 3970 14968 3976 15020
rect 4028 14968 4034 15020
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4120 14980 4646 15008
rect 4120 14968 4126 14980
rect 7742 14968 7748 15020
rect 7800 14968 7806 15020
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 2746 14912 4261 14940
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 2746 14804 2774 14912
rect 4249 14909 4261 14912
rect 4295 14909 4307 14943
rect 4249 14903 4307 14909
rect 5718 14900 5724 14952
rect 5776 14900 5782 14952
rect 5994 14900 6000 14952
rect 6052 14900 6058 14952
rect 6365 14943 6423 14949
rect 6365 14909 6377 14943
rect 6411 14909 6423 14943
rect 9876 14940 9904 15107
rect 9953 15079 10011 15085
rect 9953 15045 9965 15079
rect 9999 15076 10011 15079
rect 9999 15048 10824 15076
rect 9999 15045 10011 15048
rect 9953 15039 10011 15045
rect 10796 15020 10824 15048
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 15008 10103 15011
rect 10594 15008 10600 15020
rect 10091 14980 10600 15008
rect 10091 14977 10103 14980
rect 10045 14971 10103 14977
rect 10594 14968 10600 14980
rect 10652 14968 10658 15020
rect 10778 14968 10784 15020
rect 10836 14968 10842 15020
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 11698 15008 11704 15020
rect 11204 14980 11704 15008
rect 11204 14968 11210 14980
rect 11698 14968 11704 14980
rect 11756 15008 11762 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11756 14980 11805 15008
rect 11756 14968 11762 14980
rect 11793 14977 11805 14980
rect 11839 14977 11851 15011
rect 11793 14971 11851 14977
rect 12060 15011 12118 15017
rect 12060 14977 12072 15011
rect 12106 15008 12118 15011
rect 12360 15008 12388 15116
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 12986 15104 12992 15156
rect 13044 15144 13050 15156
rect 13173 15147 13231 15153
rect 13173 15144 13185 15147
rect 13044 15116 13185 15144
rect 13044 15104 13050 15116
rect 13173 15113 13185 15116
rect 13219 15113 13231 15147
rect 13173 15107 13231 15113
rect 15565 15147 15623 15153
rect 15565 15113 15577 15147
rect 15611 15144 15623 15147
rect 15654 15144 15660 15156
rect 15611 15116 15660 15144
rect 15611 15113 15623 15116
rect 15565 15107 15623 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 19886 15104 19892 15156
rect 19944 15104 19950 15156
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 13078 15076 13084 15088
rect 12584 15048 13084 15076
rect 12584 15036 12590 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 14452 15079 14510 15085
rect 14452 15045 14464 15079
rect 14498 15076 14510 15079
rect 14642 15076 14648 15088
rect 14498 15048 14648 15076
rect 14498 15045 14510 15048
rect 14452 15039 14510 15045
rect 14642 15036 14648 15048
rect 14700 15036 14706 15088
rect 18776 15079 18834 15085
rect 18776 15045 18788 15079
rect 18822 15076 18834 15079
rect 19058 15076 19064 15088
rect 18822 15048 19064 15076
rect 18822 15045 18834 15048
rect 18776 15039 18834 15045
rect 19058 15036 19064 15048
rect 19116 15036 19122 15088
rect 12434 15008 12440 15020
rect 12106 14980 12440 15008
rect 12106 14977 12118 14980
rect 12060 14971 12118 14977
rect 12434 14968 12440 14980
rect 12492 14968 12498 15020
rect 18138 14968 18144 15020
rect 18196 15008 18202 15020
rect 18509 15011 18567 15017
rect 18509 15008 18521 15011
rect 18196 14980 18521 15008
rect 18196 14968 18202 14980
rect 18509 14977 18521 14980
rect 18555 14977 18567 15011
rect 18509 14971 18567 14977
rect 10505 14943 10563 14949
rect 10505 14940 10517 14943
rect 9876 14912 10517 14940
rect 6365 14903 6423 14909
rect 10505 14909 10517 14912
rect 10551 14909 10563 14943
rect 10505 14903 10563 14909
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 6380 14816 6408 14903
rect 10134 14832 10140 14884
rect 10192 14872 10198 14884
rect 10229 14875 10287 14881
rect 10229 14872 10241 14875
rect 10192 14844 10241 14872
rect 10192 14832 10198 14844
rect 10229 14841 10241 14844
rect 10275 14872 10287 14875
rect 10704 14872 10732 14903
rect 14182 14900 14188 14952
rect 14240 14900 14246 14952
rect 10275 14844 10732 14872
rect 10275 14841 10287 14844
rect 10229 14835 10287 14841
rect 1820 14776 2774 14804
rect 1820 14764 1826 14776
rect 3142 14764 3148 14816
rect 3200 14764 3206 14816
rect 3510 14764 3516 14816
rect 3568 14764 3574 14816
rect 4157 14807 4215 14813
rect 4157 14773 4169 14807
rect 4203 14804 4215 14807
rect 6362 14804 6368 14816
rect 4203 14776 6368 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 7650 14764 7656 14816
rect 7708 14804 7714 14816
rect 8113 14807 8171 14813
rect 8113 14804 8125 14807
rect 7708 14776 8125 14804
rect 7708 14764 7714 14776
rect 8113 14773 8125 14776
rect 8159 14773 8171 14807
rect 8113 14767 8171 14773
rect 8938 14764 8944 14816
rect 8996 14764 9002 14816
rect 9674 14764 9680 14816
rect 9732 14764 9738 14816
rect 10042 14764 10048 14816
rect 10100 14804 10106 14816
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 10100 14776 10333 14804
rect 10100 14764 10106 14776
rect 10321 14773 10333 14776
rect 10367 14773 10379 14807
rect 10321 14767 10379 14773
rect 1104 14714 20792 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 10214 14714
rect 10266 14662 10278 14714
rect 10330 14662 10342 14714
rect 10394 14662 10406 14714
rect 10458 14662 10470 14714
rect 10522 14662 16214 14714
rect 16266 14662 16278 14714
rect 16330 14662 16342 14714
rect 16394 14662 16406 14714
rect 16458 14662 16470 14714
rect 16522 14662 20792 14714
rect 1104 14640 20792 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 1670 14600 1676 14612
rect 1627 14572 1676 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 3142 14560 3148 14612
rect 3200 14560 3206 14612
rect 3605 14603 3663 14609
rect 3605 14569 3617 14603
rect 3651 14600 3663 14603
rect 3970 14600 3976 14612
rect 3651 14572 3976 14600
rect 3651 14569 3663 14572
rect 3605 14563 3663 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 10778 14560 10784 14612
rect 10836 14560 10842 14612
rect 11425 14603 11483 14609
rect 11425 14569 11437 14603
rect 11471 14600 11483 14603
rect 12434 14600 12440 14612
rect 11471 14572 12440 14600
rect 11471 14569 11483 14572
rect 11425 14563 11483 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 17129 14603 17187 14609
rect 17129 14569 17141 14603
rect 17175 14600 17187 14603
rect 17402 14600 17408 14612
rect 17175 14572 17408 14600
rect 17175 14569 17187 14572
rect 17129 14563 17187 14569
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14464 2191 14467
rect 3160 14464 3188 14560
rect 2179 14436 3188 14464
rect 7285 14467 7343 14473
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 7285 14433 7297 14467
rect 7331 14464 7343 14467
rect 7650 14464 7656 14476
rect 7331 14436 7656 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 7926 14424 7932 14476
rect 7984 14464 7990 14476
rect 8938 14464 8944 14476
rect 7984 14436 8944 14464
rect 7984 14424 7990 14436
rect 8938 14424 8944 14436
rect 8996 14464 9002 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8996 14436 9045 14464
rect 8996 14424 9002 14436
rect 9033 14433 9045 14436
rect 9079 14464 9091 14467
rect 9079 14436 10640 14464
rect 9079 14433 9091 14436
rect 9033 14427 9091 14433
rect 10612 14408 10640 14436
rect 12802 14424 12808 14476
rect 12860 14464 12866 14476
rect 14182 14464 14188 14476
rect 12860 14436 14188 14464
rect 12860 14424 12866 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 15286 14424 15292 14476
rect 15344 14424 15350 14476
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 16724 14436 16957 14464
rect 16724 14424 16730 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 17589 14467 17647 14473
rect 17589 14464 17601 14467
rect 16945 14427 17003 14433
rect 17052 14436 17601 14464
rect 1578 14356 1584 14408
rect 1636 14356 1642 14408
rect 1762 14356 1768 14408
rect 1820 14356 1826 14408
rect 1854 14356 1860 14408
rect 1912 14356 1918 14408
rect 5810 14356 5816 14408
rect 5868 14396 5874 14408
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 5868 14368 7021 14396
rect 5868 14356 5874 14368
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 10594 14356 10600 14408
rect 10652 14356 10658 14408
rect 12526 14356 12532 14408
rect 12584 14405 12590 14408
rect 12584 14359 12596 14405
rect 15304 14396 15332 14424
rect 17052 14396 17080 14436
rect 17589 14433 17601 14436
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 17126 14405 17132 14408
rect 15304 14368 17080 14396
rect 17122 14359 17132 14405
rect 17184 14396 17190 14408
rect 17604 14396 17632 14427
rect 18138 14396 18144 14408
rect 17184 14368 17264 14396
rect 17604 14368 18144 14396
rect 12584 14356 12590 14359
rect 17126 14356 17132 14359
rect 17184 14356 17190 14368
rect 4062 14328 4068 14340
rect 3358 14300 4068 14328
rect 4062 14288 4068 14300
rect 4120 14288 4126 14340
rect 5166 14288 5172 14340
rect 5224 14328 5230 14340
rect 5224 14300 6040 14328
rect 5224 14288 5230 14300
rect 6012 14260 6040 14300
rect 6914 14288 6920 14340
rect 6972 14288 6978 14340
rect 7742 14288 7748 14340
rect 7800 14288 7806 14340
rect 9306 14288 9312 14340
rect 9364 14288 9370 14340
rect 9858 14288 9864 14340
rect 9916 14288 9922 14340
rect 15556 14331 15614 14337
rect 15556 14297 15568 14331
rect 15602 14328 15614 14331
rect 15654 14328 15660 14340
rect 15602 14300 15660 14328
rect 15602 14297 15614 14300
rect 15556 14291 15614 14297
rect 15654 14288 15660 14300
rect 15712 14328 15718 14340
rect 16853 14331 16911 14337
rect 16853 14328 16865 14331
rect 15712 14300 16865 14328
rect 15712 14288 15718 14300
rect 16853 14297 16865 14300
rect 16899 14297 16911 14331
rect 17236 14328 17264 14368
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 17834 14331 17892 14337
rect 17834 14328 17846 14331
rect 17236 14300 17846 14328
rect 16853 14291 16911 14297
rect 17834 14297 17846 14300
rect 17880 14297 17892 14331
rect 17834 14291 17892 14297
rect 7650 14260 7656 14272
rect 6012 14232 7656 14260
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 8754 14220 8760 14272
rect 8812 14220 8818 14272
rect 16666 14220 16672 14272
rect 16724 14220 16730 14272
rect 17310 14220 17316 14272
rect 17368 14220 17374 14272
rect 18966 14220 18972 14272
rect 19024 14220 19030 14272
rect 1104 14170 20792 14192
rect 1104 14118 7214 14170
rect 7266 14118 7278 14170
rect 7330 14118 7342 14170
rect 7394 14118 7406 14170
rect 7458 14118 7470 14170
rect 7522 14118 13214 14170
rect 13266 14118 13278 14170
rect 13330 14118 13342 14170
rect 13394 14118 13406 14170
rect 13458 14118 13470 14170
rect 13522 14118 19214 14170
rect 19266 14118 19278 14170
rect 19330 14118 19342 14170
rect 19394 14118 19406 14170
rect 19458 14118 19470 14170
rect 19522 14118 20792 14170
rect 1104 14096 20792 14118
rect 3237 14059 3295 14065
rect 3237 14025 3249 14059
rect 3283 14056 3295 14059
rect 3326 14056 3332 14068
rect 3283 14028 3332 14056
rect 3283 14025 3295 14028
rect 3237 14019 3295 14025
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 3970 14056 3976 14068
rect 3436 14028 3976 14056
rect 3436 13920 3464 14028
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 5537 14059 5595 14065
rect 5537 14025 5549 14059
rect 5583 14056 5595 14059
rect 5718 14056 5724 14068
rect 5583 14028 5724 14056
rect 5583 14025 5595 14028
rect 5537 14019 5595 14025
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 5810 14016 5816 14068
rect 5868 14016 5874 14068
rect 6362 14056 6368 14068
rect 5920 14028 6368 14056
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 4065 13991 4123 13997
rect 4065 13988 4077 13991
rect 3568 13960 4077 13988
rect 3568 13948 3574 13960
rect 4065 13957 4077 13960
rect 4111 13957 4123 13991
rect 4065 13951 4123 13957
rect 3697 13923 3755 13929
rect 3697 13920 3709 13923
rect 3436 13892 3709 13920
rect 3697 13889 3709 13892
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 3786 13880 3792 13932
rect 3844 13880 3850 13932
rect 5626 13920 5632 13932
rect 5198 13906 5632 13920
rect 5184 13892 5632 13906
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 5184 13852 5212 13892
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13920 5779 13923
rect 5920 13920 5948 14028
rect 6362 14016 6368 14028
rect 6420 14056 6426 14068
rect 6420 14028 7052 14056
rect 6420 14016 6426 14028
rect 6196 13960 6868 13988
rect 5767 13892 5948 13920
rect 5997 13923 6055 13929
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6086 13920 6092 13932
rect 6043 13892 6092 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 6196 13929 6224 13960
rect 6181 13923 6239 13929
rect 6181 13889 6193 13923
rect 6227 13889 6239 13923
rect 6181 13883 6239 13889
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 4120 13824 5212 13852
rect 4120 13812 4126 13824
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 6380 13852 6408 13883
rect 5408 13824 6408 13852
rect 6840 13852 6868 13960
rect 6914 13948 6920 14000
rect 6972 13948 6978 14000
rect 7024 13988 7052 14028
rect 7650 14016 7656 14068
rect 7708 14016 7714 14068
rect 7760 14028 8708 14056
rect 7760 13988 7788 14028
rect 7024 13960 7788 13988
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 8680 13997 8708 14028
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 9364 14028 9965 14056
rect 9364 14016 9370 14028
rect 9953 14025 9965 14028
rect 9999 14025 10011 14059
rect 9953 14019 10011 14025
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 11756 14028 11805 14056
rect 11756 14016 11762 14028
rect 11793 14025 11805 14028
rect 11839 14056 11851 14059
rect 12802 14056 12808 14068
rect 11839 14028 12808 14056
rect 11839 14025 11851 14028
rect 11793 14019 11851 14025
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 16574 14016 16580 14068
rect 16632 14016 16638 14068
rect 18138 14016 18144 14068
rect 18196 14016 18202 14068
rect 8573 13991 8631 13997
rect 8573 13988 8585 13991
rect 7892 13960 8585 13988
rect 7892 13948 7898 13960
rect 8573 13957 8585 13960
rect 8619 13957 8631 13991
rect 8573 13951 8631 13957
rect 8665 13991 8723 13997
rect 8665 13957 8677 13991
rect 8711 13957 8723 13991
rect 8665 13951 8723 13957
rect 9401 13991 9459 13997
rect 9401 13957 9413 13991
rect 9447 13988 9459 13991
rect 9674 13988 9680 14000
rect 9447 13960 9680 13988
rect 9447 13957 9459 13960
rect 9401 13951 9459 13957
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 14550 13948 14556 14000
rect 14608 13948 14614 14000
rect 16301 13991 16359 13997
rect 16301 13957 16313 13991
rect 16347 13988 16359 13991
rect 16592 13988 16620 14016
rect 16669 13991 16727 13997
rect 16669 13988 16681 13991
rect 16347 13960 16681 13988
rect 16347 13957 16359 13960
rect 16301 13951 16359 13957
rect 16669 13957 16681 13960
rect 16715 13957 16727 13991
rect 16669 13951 16727 13957
rect 18868 13991 18926 13997
rect 18868 13957 18880 13991
rect 18914 13988 18926 13991
rect 18966 13988 18972 14000
rect 18914 13960 18972 13988
rect 18914 13957 18926 13960
rect 18868 13951 18926 13957
rect 6932 13920 6960 13948
rect 8429 13923 8487 13929
rect 8429 13920 8441 13923
rect 6932 13892 8441 13920
rect 8429 13889 8441 13892
rect 8475 13889 8487 13923
rect 8429 13883 8487 13889
rect 8754 13880 8760 13932
rect 8812 13920 8818 13932
rect 8849 13923 8907 13929
rect 8849 13920 8861 13923
rect 8812 13892 8861 13920
rect 8812 13880 8818 13892
rect 8849 13889 8861 13892
rect 8895 13889 8907 13923
rect 8849 13883 8907 13889
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 15746 13920 15752 13932
rect 13311 13892 15752 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 8864 13852 8892 13883
rect 6840 13824 8892 13852
rect 9861 13855 9919 13861
rect 5408 13812 5414 13824
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 10152 13852 10180 13883
rect 15746 13880 15752 13892
rect 15804 13920 15810 13932
rect 16316 13920 16344 13951
rect 18966 13948 18972 13960
rect 19024 13948 19030 14000
rect 15804 13892 16344 13920
rect 15804 13880 15810 13892
rect 9907 13824 10180 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 18046 13812 18052 13864
rect 18104 13852 18110 13864
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18104 13824 18613 13852
rect 18104 13812 18110 13824
rect 18601 13821 18613 13824
rect 18647 13821 18659 13855
rect 18601 13815 18659 13821
rect 1578 13744 1584 13796
rect 1636 13784 1642 13796
rect 2682 13784 2688 13796
rect 1636 13756 2688 13784
rect 1636 13744 1642 13756
rect 2682 13744 2688 13756
rect 2740 13784 2746 13796
rect 3329 13787 3387 13793
rect 3329 13784 3341 13787
rect 2740 13756 3341 13784
rect 2740 13744 2746 13756
rect 3329 13753 3341 13756
rect 3375 13753 3387 13787
rect 3329 13747 3387 13753
rect 9769 13787 9827 13793
rect 9769 13753 9781 13787
rect 9815 13784 9827 13787
rect 10042 13784 10048 13796
rect 9815 13756 10048 13784
rect 9815 13753 9827 13756
rect 9769 13747 9827 13753
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 5994 13676 6000 13728
rect 6052 13676 6058 13728
rect 8294 13676 8300 13728
rect 8352 13676 8358 13728
rect 10505 13719 10563 13725
rect 10505 13685 10517 13719
rect 10551 13716 10563 13719
rect 10594 13716 10600 13728
rect 10551 13688 10600 13716
rect 10551 13685 10563 13688
rect 10505 13679 10563 13685
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 17126 13716 17132 13728
rect 16632 13688 17132 13716
rect 16632 13676 16638 13688
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 19978 13676 19984 13728
rect 20036 13676 20042 13728
rect 1104 13626 20792 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 10214 13626
rect 10266 13574 10278 13626
rect 10330 13574 10342 13626
rect 10394 13574 10406 13626
rect 10458 13574 10470 13626
rect 10522 13574 16214 13626
rect 16266 13574 16278 13626
rect 16330 13574 16342 13626
rect 16394 13574 16406 13626
rect 16458 13574 16470 13626
rect 16522 13574 20792 13626
rect 1104 13552 20792 13574
rect 4788 13515 4846 13521
rect 4788 13481 4800 13515
rect 4834 13512 4846 13515
rect 5994 13512 6000 13524
rect 4834 13484 6000 13512
rect 4834 13481 4846 13484
rect 4788 13475 4846 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 8113 13515 8171 13521
rect 8113 13512 8125 13515
rect 7892 13484 8125 13512
rect 7892 13472 7898 13484
rect 8113 13481 8125 13484
rect 8159 13481 8171 13515
rect 17034 13512 17040 13524
rect 8113 13475 8171 13481
rect 13004 13484 17040 13512
rect 4522 13336 4528 13388
rect 4580 13376 4586 13388
rect 5442 13376 5448 13388
rect 4580 13348 5448 13376
rect 4580 13336 4586 13348
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13376 6331 13379
rect 6641 13379 6699 13385
rect 6641 13376 6653 13379
rect 6319 13348 6653 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 6641 13345 6653 13348
rect 6687 13345 6699 13379
rect 6641 13339 6699 13345
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9732 13348 9781 13376
rect 9732 13336 9738 13348
rect 9769 13345 9781 13348
rect 9815 13376 9827 13379
rect 9950 13376 9956 13388
rect 9815 13348 9956 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10594 13376 10600 13388
rect 10367 13348 10600 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 2682 13268 2688 13320
rect 2740 13308 2746 13320
rect 3329 13311 3387 13317
rect 3329 13308 3341 13311
rect 2740 13280 3341 13308
rect 2740 13268 2746 13280
rect 3329 13277 3341 13280
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3510 13268 3516 13320
rect 3568 13268 3574 13320
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 4172 13280 4261 13308
rect 4172 13184 4200 13280
rect 4249 13277 4261 13280
rect 4295 13277 4307 13311
rect 4249 13271 4307 13277
rect 6362 13268 6368 13320
rect 6420 13268 6426 13320
rect 7742 13268 7748 13320
rect 7800 13268 7806 13320
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 9490 13308 9496 13320
rect 9171 13280 9496 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 9490 13268 9496 13280
rect 9548 13268 9554 13320
rect 9858 13268 9864 13320
rect 9916 13268 9922 13320
rect 6026 13212 6960 13240
rect 6932 13184 6960 13212
rect 2498 13132 2504 13184
rect 2556 13132 2562 13184
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 3421 13175 3479 13181
rect 3421 13172 3433 13175
rect 3200 13144 3433 13172
rect 3200 13132 3206 13144
rect 3421 13141 3433 13144
rect 3467 13141 3479 13175
rect 3421 13135 3479 13141
rect 4154 13132 4160 13184
rect 4212 13132 4218 13184
rect 4338 13132 4344 13184
rect 4396 13132 4402 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7760 13172 7788 13268
rect 9306 13200 9312 13252
rect 9364 13200 9370 13252
rect 9766 13200 9772 13252
rect 9824 13200 9830 13252
rect 10244 13240 10272 13339
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 13004 13385 13032 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17402 13472 17408 13524
rect 17460 13512 17466 13524
rect 17862 13512 17868 13524
rect 17460 13484 17868 13512
rect 17460 13472 17466 13484
rect 17862 13472 17868 13484
rect 17920 13512 17926 13524
rect 18049 13515 18107 13521
rect 18049 13512 18061 13515
rect 17920 13484 18061 13512
rect 17920 13472 17926 13484
rect 18049 13481 18061 13484
rect 18095 13481 18107 13515
rect 18049 13475 18107 13481
rect 15654 13404 15660 13456
rect 15712 13404 15718 13456
rect 16485 13447 16543 13453
rect 16485 13413 16497 13447
rect 16531 13444 16543 13447
rect 16574 13444 16580 13456
rect 16531 13416 16580 13444
rect 16531 13413 16543 13416
rect 16485 13407 16543 13413
rect 16574 13404 16580 13416
rect 16632 13404 16638 13456
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13345 13047 13379
rect 12989 13339 13047 13345
rect 14182 13336 14188 13388
rect 14240 13376 14246 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 14240 13348 14289 13376
rect 14240 13336 14246 13348
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13403 13280 15608 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 10597 13243 10655 13249
rect 10597 13240 10609 13243
rect 10244 13212 10609 13240
rect 10597 13209 10609 13212
rect 10643 13209 10655 13243
rect 10870 13240 10876 13252
rect 10597 13203 10655 13209
rect 10704 13212 10876 13240
rect 6972 13144 7788 13172
rect 6972 13132 6978 13144
rect 8938 13132 8944 13184
rect 8996 13132 9002 13184
rect 9784 13172 9812 13200
rect 10704 13172 10732 13212
rect 10870 13200 10876 13212
rect 10928 13240 10934 13252
rect 10928 13212 11086 13240
rect 10928 13200 10934 13212
rect 12158 13200 12164 13252
rect 12216 13200 12222 13252
rect 14550 13249 14556 13252
rect 13909 13243 13967 13249
rect 13909 13209 13921 13243
rect 13955 13240 13967 13243
rect 14533 13243 14556 13249
rect 14533 13240 14545 13243
rect 13955 13212 14545 13240
rect 13955 13209 13967 13212
rect 13909 13203 13967 13209
rect 14533 13209 14545 13212
rect 14533 13203 14556 13209
rect 14550 13200 14556 13203
rect 14608 13200 14614 13252
rect 9784 13144 10732 13172
rect 12066 13132 12072 13184
rect 12124 13132 12130 13184
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 13136 13144 13553 13172
rect 13136 13132 13142 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 13541 13135 13599 13141
rect 13630 13132 13636 13184
rect 13688 13132 13694 13184
rect 13722 13132 13728 13184
rect 13780 13132 13786 13184
rect 15580 13172 15608 13280
rect 15672 13240 15700 13404
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16574 13308 16580 13320
rect 15979 13280 16580 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 16669 13311 16727 13317
rect 16669 13277 16681 13311
rect 16715 13308 16727 13311
rect 17678 13308 17684 13320
rect 16715 13280 17684 13308
rect 16715 13277 16727 13280
rect 16669 13271 16727 13277
rect 17678 13268 17684 13280
rect 17736 13308 17742 13320
rect 18046 13308 18052 13320
rect 17736 13280 18052 13308
rect 17736 13268 17742 13280
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 16117 13243 16175 13249
rect 16117 13240 16129 13243
rect 15672 13212 16129 13240
rect 16117 13209 16129 13212
rect 16163 13209 16175 13243
rect 16117 13203 16175 13209
rect 16209 13243 16267 13249
rect 16209 13209 16221 13243
rect 16255 13240 16267 13243
rect 16914 13243 16972 13249
rect 16914 13240 16926 13243
rect 16255 13212 16436 13240
rect 16255 13209 16267 13212
rect 16209 13203 16267 13209
rect 16022 13172 16028 13184
rect 15580 13144 16028 13172
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 16298 13132 16304 13184
rect 16356 13132 16362 13184
rect 16408 13172 16436 13212
rect 16776 13212 16926 13240
rect 16666 13172 16672 13184
rect 16408 13144 16672 13172
rect 16666 13132 16672 13144
rect 16724 13172 16730 13184
rect 16776 13172 16804 13212
rect 16914 13209 16926 13212
rect 16960 13209 16972 13243
rect 16914 13203 16972 13209
rect 16724 13144 16804 13172
rect 16724 13132 16730 13144
rect 1104 13082 20792 13104
rect 1104 13030 7214 13082
rect 7266 13030 7278 13082
rect 7330 13030 7342 13082
rect 7394 13030 7406 13082
rect 7458 13030 7470 13082
rect 7522 13030 13214 13082
rect 13266 13030 13278 13082
rect 13330 13030 13342 13082
rect 13394 13030 13406 13082
rect 13458 13030 13470 13082
rect 13522 13030 19214 13082
rect 19266 13030 19278 13082
rect 19330 13030 19342 13082
rect 19394 13030 19406 13082
rect 19458 13030 19470 13082
rect 19522 13030 20792 13082
rect 1104 13008 20792 13030
rect 2682 12928 2688 12980
rect 2740 12928 2746 12980
rect 3142 12928 3148 12980
rect 3200 12928 3206 12980
rect 4338 12928 4344 12980
rect 4396 12928 4402 12980
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 7009 12971 7067 12977
rect 7009 12968 7021 12971
rect 6420 12940 7021 12968
rect 6420 12928 6426 12940
rect 7009 12937 7021 12940
rect 7055 12937 7067 12971
rect 7009 12931 7067 12937
rect 7926 12928 7932 12980
rect 7984 12928 7990 12980
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9180 12940 9781 12968
rect 9180 12928 9186 12940
rect 9769 12937 9781 12940
rect 9815 12937 9827 12971
rect 9769 12931 9827 12937
rect 2700 12900 2728 12928
rect 2148 12872 2728 12900
rect 2869 12903 2927 12909
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 1394 12724 1400 12776
rect 1452 12764 1458 12776
rect 1688 12764 1716 12795
rect 1452 12736 1716 12764
rect 1452 12724 1458 12736
rect 1670 12656 1676 12708
rect 1728 12696 1734 12708
rect 2148 12705 2176 12872
rect 2869 12869 2881 12903
rect 2915 12900 2927 12903
rect 3160 12900 3188 12928
rect 2915 12872 3188 12900
rect 2915 12869 2927 12872
rect 2869 12863 2927 12869
rect 2498 12792 2504 12844
rect 2556 12832 2562 12844
rect 2593 12835 2651 12841
rect 2593 12832 2605 12835
rect 2556 12804 2605 12832
rect 2556 12792 2562 12804
rect 2593 12801 2605 12804
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 4356 12832 4384 12928
rect 7098 12900 7104 12912
rect 6748 12872 7104 12900
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 4356 12804 4445 12832
rect 4433 12801 4445 12804
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 6748 12841 6776 12872
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 5776 12804 6377 12832
rect 5776 12792 5782 12804
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6733 12835 6791 12841
rect 6733 12801 6745 12835
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 6917 12835 6975 12841
rect 6917 12801 6929 12835
rect 6963 12801 6975 12835
rect 7944 12832 7972 12928
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7944 12804 8033 12832
rect 6917 12795 6975 12801
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 2409 12767 2467 12773
rect 2409 12733 2421 12767
rect 2455 12733 2467 12767
rect 2409 12727 2467 12733
rect 2133 12699 2191 12705
rect 2133 12696 2145 12699
rect 1728 12668 2145 12696
rect 1728 12656 1734 12668
rect 2133 12665 2145 12668
rect 2179 12665 2191 12699
rect 2133 12659 2191 12665
rect 1762 12588 1768 12640
rect 1820 12588 1826 12640
rect 1946 12588 1952 12640
rect 2004 12588 2010 12640
rect 2424 12628 2452 12727
rect 3418 12724 3424 12776
rect 3476 12764 3482 12776
rect 3988 12764 4016 12792
rect 3476 12736 4016 12764
rect 4341 12767 4399 12773
rect 3476 12724 3482 12736
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4709 12767 4767 12773
rect 4709 12764 4721 12767
rect 4387 12736 4721 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 4709 12733 4721 12736
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 6932 12764 6960 12795
rect 9398 12792 9404 12844
rect 9456 12832 9462 12844
rect 9784 12832 9812 12931
rect 9858 12928 9864 12980
rect 9916 12968 9922 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 9916 12940 10701 12968
rect 9916 12928 9922 12940
rect 10689 12937 10701 12940
rect 10735 12937 10747 12971
rect 10689 12931 10747 12937
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 11609 12971 11667 12977
rect 11609 12968 11621 12971
rect 10928 12940 11621 12968
rect 10928 12928 10934 12940
rect 11609 12937 11621 12940
rect 11655 12937 11667 12971
rect 11609 12931 11667 12937
rect 12066 12928 12072 12980
rect 12124 12928 12130 12980
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 13630 12968 13636 12980
rect 12299 12940 13636 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 13630 12928 13636 12940
rect 13688 12968 13694 12980
rect 14090 12968 14096 12980
rect 13688 12940 14096 12968
rect 13688 12928 13694 12940
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 14550 12968 14556 12980
rect 14231 12940 14556 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 14550 12928 14556 12940
rect 14608 12968 14614 12980
rect 14608 12940 15792 12968
rect 14608 12928 14614 12940
rect 9950 12860 9956 12912
rect 10008 12900 10014 12912
rect 10137 12903 10195 12909
rect 10137 12900 10149 12903
rect 10008 12872 10149 12900
rect 10008 12860 10014 12872
rect 10137 12869 10149 12872
rect 10183 12869 10195 12903
rect 12084 12900 12112 12928
rect 15286 12900 15292 12912
rect 15344 12909 15350 12912
rect 10137 12863 10195 12869
rect 11348 12872 12112 12900
rect 15256 12872 15292 12900
rect 11348 12841 11376 12872
rect 15286 12860 15292 12872
rect 15344 12863 15356 12909
rect 15396 12872 15700 12900
rect 15344 12860 15350 12863
rect 10505 12835 10563 12841
rect 10505 12832 10517 12835
rect 9456 12804 9628 12832
rect 9784 12804 10517 12832
rect 9456 12792 9462 12804
rect 5500 12736 6960 12764
rect 8297 12767 8355 12773
rect 5500 12724 5506 12736
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 8386 12764 8392 12776
rect 8343 12736 8392 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 9490 12724 9496 12776
rect 9548 12724 9554 12776
rect 9600 12764 9628 12804
rect 10505 12801 10517 12804
rect 10551 12801 10563 12835
rect 10505 12795 10563 12801
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 9766 12764 9772 12776
rect 9600 12736 9772 12764
rect 9766 12724 9772 12736
rect 9824 12724 9830 12776
rect 9508 12696 9536 12724
rect 9953 12699 10011 12705
rect 9953 12696 9965 12699
rect 9508 12668 9965 12696
rect 9953 12665 9965 12668
rect 9999 12665 10011 12699
rect 9953 12659 10011 12665
rect 4706 12628 4712 12640
rect 2424 12600 4712 12628
rect 4706 12588 4712 12600
rect 4764 12628 4770 12640
rect 6181 12631 6239 12637
rect 6181 12628 6193 12631
rect 4764 12600 6193 12628
rect 4764 12588 4770 12600
rect 6181 12597 6193 12600
rect 6227 12597 6239 12631
rect 6181 12591 6239 12597
rect 10134 12588 10140 12640
rect 10192 12628 10198 12640
rect 11348 12628 11376 12795
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13366 12835 13424 12841
rect 13366 12832 13378 12835
rect 13136 12804 13378 12832
rect 13136 12792 13142 12804
rect 13366 12801 13378 12804
rect 13412 12832 13424 12835
rect 15396 12832 15424 12872
rect 15672 12841 15700 12872
rect 13412 12804 15424 12832
rect 15657 12835 15715 12841
rect 13412 12801 13424 12804
rect 13366 12795 13424 12801
rect 15657 12801 15669 12835
rect 15703 12801 15715 12835
rect 15764 12832 15792 12940
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 16666 12968 16672 12980
rect 16080 12940 16672 12968
rect 16080 12928 16086 12940
rect 16666 12928 16672 12940
rect 16724 12928 16730 12980
rect 16761 12971 16819 12977
rect 16761 12937 16773 12971
rect 16807 12968 16819 12971
rect 17126 12968 17132 12980
rect 16807 12940 17132 12968
rect 16807 12937 16819 12940
rect 16761 12931 16819 12937
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 18693 12971 18751 12977
rect 18693 12937 18705 12971
rect 18739 12968 18751 12971
rect 19242 12968 19248 12980
rect 18739 12940 19248 12968
rect 18739 12937 18751 12940
rect 18693 12931 18751 12937
rect 19242 12928 19248 12940
rect 19300 12968 19306 12980
rect 20349 12971 20407 12977
rect 20349 12968 20361 12971
rect 19300 12940 20361 12968
rect 19300 12928 19306 12940
rect 20349 12937 20361 12940
rect 20395 12937 20407 12971
rect 20349 12931 20407 12937
rect 16298 12860 16304 12912
rect 16356 12900 16362 12912
rect 17862 12900 17868 12912
rect 17920 12909 17926 12912
rect 16356 12872 17868 12900
rect 16356 12860 16362 12872
rect 17862 12860 17868 12872
rect 17920 12900 17932 12909
rect 17920 12872 17965 12900
rect 17920 12863 17932 12872
rect 17920 12860 17926 12863
rect 18506 12860 18512 12912
rect 18564 12900 18570 12912
rect 18966 12900 18972 12912
rect 18564 12872 18972 12900
rect 18564 12860 18570 12872
rect 18966 12860 18972 12872
rect 19024 12860 19030 12912
rect 19978 12860 19984 12912
rect 20036 12860 20042 12912
rect 15933 12835 15991 12841
rect 15933 12832 15945 12835
rect 15764 12804 15945 12832
rect 15657 12795 15715 12801
rect 15933 12801 15945 12804
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 18046 12792 18052 12844
rect 18104 12832 18110 12844
rect 18141 12835 18199 12841
rect 18141 12832 18153 12835
rect 18104 12804 18153 12832
rect 18104 12792 18110 12804
rect 18141 12801 18153 12804
rect 18187 12801 18199 12835
rect 18141 12795 18199 12801
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12832 18659 12835
rect 19236 12835 19294 12841
rect 19236 12832 19248 12835
rect 18647 12804 19248 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 19236 12801 19248 12804
rect 19282 12832 19294 12835
rect 19518 12832 19524 12844
rect 19282 12804 19524 12832
rect 19282 12801 19294 12804
rect 19236 12795 19294 12801
rect 13630 12724 13636 12776
rect 13688 12724 13694 12776
rect 15562 12724 15568 12776
rect 15620 12724 15626 12776
rect 15841 12767 15899 12773
rect 15841 12764 15853 12767
rect 15672 12736 15853 12764
rect 15672 12708 15700 12736
rect 15841 12733 15853 12736
rect 15887 12733 15899 12767
rect 18156 12764 18184 12795
rect 19518 12792 19524 12804
rect 19576 12832 19582 12844
rect 19996 12832 20024 12860
rect 19576 12804 20024 12832
rect 19576 12792 19582 12804
rect 18782 12764 18788 12776
rect 18156 12736 18788 12764
rect 15841 12727 15899 12733
rect 18782 12724 18788 12736
rect 18840 12764 18846 12776
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 18840 12736 18981 12764
rect 18840 12724 18846 12736
rect 18969 12733 18981 12736
rect 19015 12733 19027 12767
rect 18969 12727 19027 12733
rect 15654 12656 15660 12708
rect 15712 12656 15718 12708
rect 17126 12696 17132 12708
rect 16132 12668 17132 12696
rect 10192 12600 11376 12628
rect 10192 12588 10198 12600
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 15286 12628 15292 12640
rect 13780 12600 15292 12628
rect 13780 12588 13786 12600
rect 15286 12588 15292 12600
rect 15344 12628 15350 12640
rect 16132 12637 16160 12668
rect 17126 12656 17132 12668
rect 17184 12656 17190 12708
rect 18874 12656 18880 12708
rect 18932 12656 18938 12708
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15344 12600 15761 12628
rect 15344 12588 15350 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 16117 12631 16175 12637
rect 16117 12597 16129 12631
rect 16163 12597 16175 12631
rect 16117 12591 16175 12597
rect 18322 12588 18328 12640
rect 18380 12588 18386 12640
rect 1104 12538 20792 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 10214 12538
rect 10266 12486 10278 12538
rect 10330 12486 10342 12538
rect 10394 12486 10406 12538
rect 10458 12486 10470 12538
rect 10522 12486 16214 12538
rect 16266 12486 16278 12538
rect 16330 12486 16342 12538
rect 16394 12486 16406 12538
rect 16458 12486 16470 12538
rect 16522 12486 20792 12538
rect 1104 12464 20792 12486
rect 1946 12384 1952 12436
rect 2004 12384 2010 12436
rect 3510 12384 3516 12436
rect 3568 12424 3574 12436
rect 3605 12427 3663 12433
rect 3605 12424 3617 12427
rect 3568 12396 3617 12424
rect 3568 12384 3574 12396
rect 3605 12393 3617 12396
rect 3651 12393 3663 12427
rect 3605 12387 3663 12393
rect 4341 12427 4399 12433
rect 4341 12393 4353 12427
rect 4387 12424 4399 12427
rect 5350 12424 5356 12436
rect 4387 12396 5356 12424
rect 4387 12393 4399 12396
rect 4341 12387 4399 12393
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8444 12396 8585 12424
rect 8444 12384 8450 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 9306 12384 9312 12436
rect 9364 12384 9370 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14185 12427 14243 12433
rect 14185 12424 14197 12427
rect 13780 12396 14197 12424
rect 13780 12384 13786 12396
rect 14185 12393 14197 12396
rect 14231 12393 14243 12427
rect 14185 12387 14243 12393
rect 19242 12384 19248 12436
rect 19300 12384 19306 12436
rect 20073 12427 20131 12433
rect 20073 12424 20085 12427
rect 19352 12396 20085 12424
rect 1964 12288 1992 12384
rect 18598 12316 18604 12368
rect 18656 12356 18662 12368
rect 18969 12359 19027 12365
rect 18969 12356 18981 12359
rect 18656 12328 18981 12356
rect 18656 12316 18662 12328
rect 18969 12325 18981 12328
rect 19015 12356 19027 12359
rect 19352 12356 19380 12396
rect 20073 12393 20085 12396
rect 20119 12393 20131 12427
rect 20073 12387 20131 12393
rect 19015 12328 19380 12356
rect 19015 12325 19027 12328
rect 18969 12319 19027 12325
rect 19518 12316 19524 12368
rect 19576 12316 19582 12368
rect 19705 12359 19763 12365
rect 19705 12325 19717 12359
rect 19751 12356 19763 12359
rect 19981 12359 20039 12365
rect 19981 12356 19993 12359
rect 19751 12328 19993 12356
rect 19751 12325 19763 12328
rect 19705 12319 19763 12325
rect 19981 12325 19993 12328
rect 20027 12325 20039 12359
rect 19981 12319 20039 12325
rect 1780 12260 1992 12288
rect 1394 12180 1400 12232
rect 1452 12180 1458 12232
rect 1780 12229 1808 12260
rect 2590 12248 2596 12300
rect 2648 12288 2654 12300
rect 2648 12260 4108 12288
rect 2648 12248 2654 12260
rect 1765 12223 1823 12229
rect 1765 12189 1777 12223
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 1854 12180 1860 12232
rect 1912 12180 1918 12232
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3789 12223 3847 12229
rect 3789 12220 3801 12223
rect 3436 12192 3801 12220
rect 1412 12152 1440 12180
rect 2133 12155 2191 12161
rect 1412 12124 2084 12152
rect 1578 12044 1584 12096
rect 1636 12044 1642 12096
rect 2056 12084 2084 12124
rect 2133 12121 2145 12155
rect 2179 12152 2191 12155
rect 2406 12152 2412 12164
rect 2179 12124 2412 12152
rect 2179 12121 2191 12124
rect 2133 12115 2191 12121
rect 2406 12112 2412 12124
rect 2464 12112 2470 12164
rect 3436 12084 3464 12192
rect 3789 12189 3801 12192
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 4080 12164 4108 12260
rect 17586 12248 17592 12300
rect 17644 12248 17650 12300
rect 18874 12288 18880 12300
rect 18616 12260 18880 12288
rect 4209 12223 4267 12229
rect 4209 12189 4221 12223
rect 4255 12220 4267 12223
rect 4706 12220 4712 12232
rect 4255 12192 4712 12220
rect 4255 12189 4267 12192
rect 4209 12183 4267 12189
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 8754 12180 8760 12232
rect 8812 12180 8818 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9582 12180 9588 12232
rect 9640 12180 9646 12232
rect 10134 12180 10140 12232
rect 10192 12180 10198 12232
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 12768 12192 13277 12220
rect 12768 12180 12774 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 14090 12180 14096 12232
rect 14148 12180 14154 12232
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 15562 12220 15568 12232
rect 14424 12192 15568 12220
rect 14424 12180 14430 12192
rect 15562 12180 15568 12192
rect 15620 12220 15626 12232
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15620 12192 15669 12220
rect 15620 12180 15626 12192
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 17856 12223 17914 12229
rect 17856 12189 17868 12223
rect 17902 12220 17914 12223
rect 18616 12220 18644 12260
rect 18874 12248 18880 12260
rect 18932 12288 18938 12300
rect 19429 12291 19487 12297
rect 18932 12260 19380 12288
rect 18932 12248 18938 12260
rect 17902 12192 18644 12220
rect 17902 12189 17914 12192
rect 17856 12183 17914 12189
rect 18690 12180 18696 12232
rect 18748 12220 18754 12232
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 18748 12192 19257 12220
rect 18748 12180 18754 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19352 12220 19380 12260
rect 19429 12257 19441 12291
rect 19475 12288 19487 12291
rect 19536 12288 19564 12316
rect 19475 12260 19564 12288
rect 19475 12257 19487 12260
rect 19429 12251 19487 12257
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 19352 12192 19533 12220
rect 19245 12183 19303 12189
rect 19521 12189 19533 12192
rect 19567 12220 19579 12223
rect 19567 12192 20852 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 3510 12112 3516 12164
rect 3568 12152 3574 12164
rect 3973 12155 4031 12161
rect 3973 12152 3985 12155
rect 3568 12124 3985 12152
rect 3568 12112 3574 12124
rect 3973 12121 3985 12124
rect 4019 12121 4031 12155
rect 3973 12115 4031 12121
rect 4062 12112 4068 12164
rect 4120 12152 4126 12164
rect 5258 12152 5264 12164
rect 4120 12124 5264 12152
rect 4120 12112 4126 12124
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 9493 12155 9551 12161
rect 9493 12121 9505 12155
rect 9539 12152 9551 12155
rect 10152 12152 10180 12180
rect 9539 12124 10180 12152
rect 14108 12152 14136 12180
rect 15930 12161 15936 12164
rect 15298 12155 15356 12161
rect 15298 12152 15310 12155
rect 14108 12124 15310 12152
rect 9539 12121 9551 12124
rect 9493 12115 9551 12121
rect 15298 12121 15310 12124
rect 15344 12121 15356 12155
rect 15924 12152 15936 12161
rect 15891 12124 15936 12152
rect 15298 12115 15356 12121
rect 15924 12115 15936 12124
rect 2056 12056 3464 12084
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12713 12087 12771 12093
rect 12713 12084 12725 12087
rect 12584 12056 12725 12084
rect 12584 12044 12590 12056
rect 12713 12053 12725 12056
rect 12759 12053 12771 12087
rect 15313 12084 15341 12115
rect 15930 12112 15936 12115
rect 15988 12112 15994 12164
rect 18046 12112 18052 12164
rect 18104 12152 18110 12164
rect 19797 12155 19855 12161
rect 19797 12152 19809 12155
rect 18104 12124 19809 12152
rect 18104 12112 18110 12124
rect 19797 12121 19809 12124
rect 19843 12121 19855 12155
rect 19797 12115 19855 12121
rect 20162 12112 20168 12164
rect 20220 12112 20226 12164
rect 15654 12084 15660 12096
rect 15313 12056 15660 12084
rect 12713 12047 12771 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16666 12044 16672 12096
rect 16724 12084 16730 12096
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 16724 12056 17049 12084
rect 16724 12044 16730 12056
rect 17037 12053 17049 12056
rect 17083 12084 17095 12087
rect 18138 12084 18144 12096
rect 17083 12056 18144 12084
rect 17083 12053 17095 12056
rect 17037 12047 17095 12053
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 19886 12044 19892 12096
rect 19944 12044 19950 12096
rect 1104 11994 20792 12016
rect 1104 11942 7214 11994
rect 7266 11942 7278 11994
rect 7330 11942 7342 11994
rect 7394 11942 7406 11994
rect 7458 11942 7470 11994
rect 7522 11942 13214 11994
rect 13266 11942 13278 11994
rect 13330 11942 13342 11994
rect 13394 11942 13406 11994
rect 13458 11942 13470 11994
rect 13522 11942 19214 11994
rect 19266 11942 19278 11994
rect 19330 11942 19342 11994
rect 19394 11942 19406 11994
rect 19458 11942 19470 11994
rect 19522 11942 20792 11994
rect 1104 11920 20792 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 1636 11852 1716 11880
rect 1636 11840 1642 11852
rect 1688 11821 1716 11852
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 2464 11852 3157 11880
rect 2464 11840 2470 11852
rect 3145 11849 3157 11852
rect 3191 11849 3203 11883
rect 3145 11843 3203 11849
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 4062 11880 4068 11892
rect 3743 11852 4068 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 13078 11880 13084 11892
rect 12207 11852 13084 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 13630 11840 13636 11892
rect 13688 11840 13694 11892
rect 16209 11883 16267 11889
rect 16209 11849 16221 11883
rect 16255 11880 16267 11883
rect 16255 11852 16712 11880
rect 16255 11849 16267 11852
rect 16209 11843 16267 11849
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11781 1731 11815
rect 13648 11812 13676 11840
rect 14366 11812 14372 11824
rect 1673 11775 1731 11781
rect 13556 11784 14372 11812
rect 1394 11704 1400 11756
rect 1452 11704 1458 11756
rect 3418 11744 3424 11756
rect 2806 11716 3424 11744
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 8662 11704 8668 11756
rect 8720 11704 8726 11756
rect 9766 11704 9772 11756
rect 9824 11704 9830 11756
rect 13556 11753 13584 11784
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 15841 11815 15899 11821
rect 15841 11781 15853 11815
rect 15887 11781 15899 11815
rect 15841 11775 15899 11781
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11713 11115 11747
rect 11057 11707 11115 11713
rect 13285 11747 13343 11753
rect 13285 11713 13297 11747
rect 13331 11744 13343 11747
rect 13541 11747 13599 11753
rect 13331 11716 13492 11744
rect 13331 11713 13343 11716
rect 13285 11707 13343 11713
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 8938 11676 8944 11688
rect 6880 11648 8944 11676
rect 6880 11636 6886 11648
rect 8938 11636 8944 11648
rect 8996 11676 9002 11688
rect 11072 11676 11100 11707
rect 11146 11676 11152 11688
rect 8996 11648 11152 11676
rect 8996 11636 9002 11648
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 13464 11676 13492 11716
rect 13541 11713 13553 11747
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11744 13691 11747
rect 15746 11744 15752 11756
rect 13679 11716 15752 11744
rect 13679 11713 13691 11716
rect 13633 11707 13691 11713
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 15856 11676 15884 11775
rect 15930 11772 15936 11824
rect 15988 11812 15994 11824
rect 16684 11821 16712 11852
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 16869 11883 16927 11889
rect 16869 11880 16881 11883
rect 16816 11852 16881 11880
rect 16816 11840 16822 11852
rect 16869 11849 16881 11852
rect 16915 11849 16927 11883
rect 16869 11843 16927 11849
rect 17497 11883 17555 11889
rect 17497 11849 17509 11883
rect 17543 11880 17555 11883
rect 18046 11880 18052 11892
rect 17543 11852 18052 11880
rect 17543 11849 17555 11852
rect 17497 11843 17555 11849
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 19886 11880 19892 11892
rect 18156 11852 19892 11880
rect 16041 11815 16099 11821
rect 16041 11812 16053 11815
rect 15988 11784 16053 11812
rect 15988 11772 15994 11784
rect 16041 11781 16053 11784
rect 16087 11781 16099 11815
rect 16041 11775 16099 11781
rect 16669 11815 16727 11821
rect 16669 11781 16681 11815
rect 16715 11781 16727 11815
rect 16669 11775 16727 11781
rect 17954 11772 17960 11824
rect 18012 11772 18018 11824
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 17310 11744 17316 11756
rect 17175 11716 17316 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 18156 11753 18184 11852
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 20349 11883 20407 11889
rect 20349 11849 20361 11883
rect 20395 11880 20407 11883
rect 20824 11880 20852 12192
rect 20395 11852 20852 11880
rect 20395 11849 20407 11852
rect 20349 11843 20407 11849
rect 18509 11815 18567 11821
rect 18509 11781 18521 11815
rect 18555 11812 18567 11815
rect 18598 11812 18604 11824
rect 18555 11784 18604 11812
rect 18555 11781 18567 11784
rect 18509 11775 18567 11781
rect 18598 11772 18604 11784
rect 18656 11772 18662 11824
rect 19058 11772 19064 11824
rect 19116 11812 19122 11824
rect 19214 11815 19272 11821
rect 19214 11812 19226 11815
rect 19116 11784 19226 11812
rect 19116 11772 19122 11784
rect 19214 11781 19226 11784
rect 19260 11781 19272 11815
rect 19214 11775 19272 11781
rect 20162 11772 20168 11824
rect 20220 11772 20226 11824
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 18322 11704 18328 11756
rect 18380 11704 18386 11756
rect 18966 11704 18972 11756
rect 19024 11704 19030 11756
rect 20180 11744 20208 11772
rect 19076 11716 20208 11744
rect 13464 11648 15884 11676
rect 15856 11608 15884 11648
rect 17218 11636 17224 11688
rect 17276 11636 17282 11688
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11645 18291 11679
rect 18340 11676 18368 11704
rect 18417 11679 18475 11685
rect 18417 11676 18429 11679
rect 18340 11648 18429 11676
rect 18233 11639 18291 11645
rect 18417 11645 18429 11648
rect 18463 11645 18475 11679
rect 18417 11639 18475 11645
rect 18601 11679 18659 11685
rect 18601 11645 18613 11679
rect 18647 11676 18659 11679
rect 19076 11676 19104 11716
rect 18647 11648 19104 11676
rect 18647 11645 18659 11648
rect 18601 11639 18659 11645
rect 16758 11608 16764 11620
rect 15856 11580 16764 11608
rect 16758 11568 16764 11580
rect 16816 11568 16822 11620
rect 17037 11611 17095 11617
rect 17037 11577 17049 11611
rect 17083 11608 17095 11611
rect 18248 11608 18276 11639
rect 17083 11580 18276 11608
rect 17083 11577 17095 11580
rect 17037 11571 17095 11577
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 8481 11543 8539 11549
rect 8481 11540 8493 11543
rect 8444 11512 8493 11540
rect 8444 11500 8450 11512
rect 8481 11509 8493 11512
rect 8527 11509 8539 11543
rect 8481 11503 8539 11509
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9916 11512 9965 11540
rect 9916 11500 9922 11512
rect 9953 11509 9965 11512
rect 9999 11509 10011 11543
rect 9953 11503 10011 11509
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 10965 11543 11023 11549
rect 10965 11540 10977 11543
rect 10928 11512 10977 11540
rect 10928 11500 10934 11512
rect 10965 11509 10977 11512
rect 11011 11509 11023 11543
rect 10965 11503 11023 11509
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14921 11543 14979 11549
rect 14921 11540 14933 11543
rect 14424 11512 14933 11540
rect 14424 11500 14430 11512
rect 14921 11509 14933 11512
rect 14967 11509 14979 11543
rect 14921 11503 14979 11509
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 16666 11540 16672 11552
rect 16071 11512 16672 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16850 11500 16856 11552
rect 16908 11500 16914 11552
rect 17126 11500 17132 11552
rect 17184 11500 17190 11552
rect 1104 11450 20792 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 10214 11450
rect 10266 11398 10278 11450
rect 10330 11398 10342 11450
rect 10394 11398 10406 11450
rect 10458 11398 10470 11450
rect 10522 11398 16214 11450
rect 16266 11398 16278 11450
rect 16330 11398 16342 11450
rect 16394 11398 16406 11450
rect 16458 11398 16470 11450
rect 16522 11398 20792 11450
rect 1104 11376 20792 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1670 11336 1676 11348
rect 1627 11308 1676 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 5169 11339 5227 11345
rect 5169 11305 5181 11339
rect 5215 11336 5227 11339
rect 5258 11336 5264 11348
rect 5215 11308 5264 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 5258 11296 5264 11308
rect 5316 11336 5322 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 5316 11308 7665 11336
rect 5316 11296 5322 11308
rect 7653 11305 7665 11308
rect 7699 11336 7711 11339
rect 7926 11336 7932 11348
rect 7699 11308 7932 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 7926 11296 7932 11308
rect 7984 11296 7990 11348
rect 8573 11339 8631 11345
rect 8573 11305 8585 11339
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 9766 11336 9772 11348
rect 8803 11308 9772 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 8588 11268 8616 11299
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 12710 11296 12716 11348
rect 12768 11296 12774 11348
rect 17218 11296 17224 11348
rect 17276 11296 17282 11348
rect 17586 11296 17592 11348
rect 17644 11336 17650 11348
rect 18046 11336 18052 11348
rect 17644 11308 18052 11336
rect 17644 11296 17650 11308
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 18138 11296 18144 11348
rect 18196 11296 18202 11348
rect 19610 11296 19616 11348
rect 19668 11296 19674 11348
rect 9030 11268 9036 11280
rect 8588 11240 9036 11268
rect 9030 11228 9036 11240
rect 9088 11228 9094 11280
rect 17236 11268 17264 11296
rect 18509 11271 18567 11277
rect 18509 11268 18521 11271
rect 17236 11240 18521 11268
rect 18509 11237 18521 11240
rect 18555 11237 18567 11271
rect 18509 11231 18567 11237
rect 19245 11271 19303 11277
rect 19245 11237 19257 11271
rect 19291 11237 19303 11271
rect 19245 11231 19303 11237
rect 5258 11160 5264 11212
rect 5316 11160 5322 11212
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9309 11203 9367 11209
rect 8996 11172 9076 11200
rect 8996 11160 9002 11172
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 6914 11132 6920 11144
rect 6670 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11132 6978 11144
rect 9048 11141 9076 11172
rect 9309 11169 9321 11203
rect 9355 11200 9367 11203
rect 10594 11200 10600 11212
rect 9355 11172 10600 11200
rect 9355 11169 9367 11172
rect 9309 11163 9367 11169
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 10781 11203 10839 11209
rect 10781 11169 10793 11203
rect 10827 11200 10839 11203
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 10827 11172 11161 11200
rect 10827 11169 10839 11172
rect 10781 11163 10839 11169
rect 11149 11169 11161 11172
rect 11195 11169 11207 11203
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 11149 11163 11207 11169
rect 12268 11172 13369 11200
rect 9033 11135 9091 11141
rect 6972 11104 7144 11132
rect 6972 11092 6978 11104
rect 5534 11024 5540 11076
rect 5592 11024 5598 11076
rect 7006 10956 7012 11008
rect 7064 10956 7070 11008
rect 7116 10996 7144 11104
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 10870 11092 10876 11144
rect 10928 11092 10934 11144
rect 8202 11024 8208 11076
rect 8260 11024 8266 11076
rect 8389 11067 8447 11073
rect 8389 11033 8401 11067
rect 8435 11064 8447 11067
rect 8478 11064 8484 11076
rect 8435 11036 8484 11064
rect 8435 11033 8447 11036
rect 8389 11027 8447 11033
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 8605 11067 8663 11073
rect 8605 11033 8617 11067
rect 8651 11064 8663 11067
rect 9398 11064 9404 11076
rect 8651 11036 9404 11064
rect 8651 11033 8663 11036
rect 8605 11027 8663 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 11054 11064 11060 11076
rect 10534 11036 11060 11064
rect 11054 11024 11060 11036
rect 11112 11064 11118 11076
rect 11112 11036 11638 11064
rect 11112 11024 11118 11036
rect 8110 10996 8116 11008
rect 7116 10968 8116 10996
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 11532 10996 11560 11036
rect 12268 10996 12296 11172
rect 13357 11169 13369 11172
rect 13403 11200 13415 11203
rect 13906 11200 13912 11212
rect 13403 11172 13912 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 19260 11200 19288 11231
rect 17828 11172 19288 11200
rect 19444 11172 19840 11200
rect 17828 11160 17834 11172
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11132 13691 11135
rect 15657 11135 15715 11141
rect 15657 11132 15669 11135
rect 13679 11104 15669 11132
rect 13679 11101 13691 11104
rect 13633 11095 13691 11101
rect 15657 11101 15669 11104
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 15930 11092 15936 11144
rect 15988 11132 15994 11144
rect 19444 11141 19472 11172
rect 19812 11144 19840 11172
rect 18141 11135 18199 11141
rect 18141 11132 18153 11135
rect 15988 11104 18153 11132
rect 15988 11092 15994 11104
rect 18141 11101 18153 11104
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 13541 11067 13599 11073
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 13814 11064 13820 11076
rect 13587 11036 13820 11064
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14093 11067 14151 11073
rect 14093 11033 14105 11067
rect 14139 11033 14151 11067
rect 14093 11027 14151 11033
rect 11532 10968 12296 10996
rect 12618 10956 12624 11008
rect 12676 10956 12682 11008
rect 13078 10956 13084 11008
rect 13136 10996 13142 11008
rect 14108 10996 14136 11027
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 16301 11067 16359 11073
rect 16301 11064 16313 11067
rect 15896 11036 16313 11064
rect 15896 11024 15902 11036
rect 16301 11033 16313 11036
rect 16347 11033 16359 11067
rect 16301 11027 16359 11033
rect 16758 11024 16764 11076
rect 16816 11064 16822 11076
rect 18248 11064 18276 11095
rect 16816 11036 18276 11064
rect 16816 11024 16822 11036
rect 13136 10968 14136 10996
rect 19536 10996 19564 11095
rect 19794 11092 19800 11144
rect 19852 11092 19858 11144
rect 19702 11024 19708 11076
rect 19760 11024 19766 11076
rect 20070 10996 20076 11008
rect 19536 10968 20076 10996
rect 13136 10956 13142 10968
rect 20070 10956 20076 10968
rect 20128 10956 20134 11008
rect 1104 10906 20792 10928
rect 1104 10854 7214 10906
rect 7266 10854 7278 10906
rect 7330 10854 7342 10906
rect 7394 10854 7406 10906
rect 7458 10854 7470 10906
rect 7522 10854 13214 10906
rect 13266 10854 13278 10906
rect 13330 10854 13342 10906
rect 13394 10854 13406 10906
rect 13458 10854 13470 10906
rect 13522 10854 19214 10906
rect 19266 10854 19278 10906
rect 19330 10854 19342 10906
rect 19394 10854 19406 10906
rect 19458 10854 19470 10906
rect 19522 10854 20792 10906
rect 1104 10832 20792 10854
rect 3237 10795 3295 10801
rect 3237 10761 3249 10795
rect 3283 10792 3295 10795
rect 4614 10792 4620 10804
rect 3283 10764 4620 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 4856 10764 5304 10792
rect 4856 10752 4862 10764
rect 4525 10727 4583 10733
rect 4525 10693 4537 10727
rect 4571 10724 4583 10727
rect 5166 10724 5172 10736
rect 4571 10696 5172 10724
rect 4571 10693 4583 10696
rect 4525 10687 4583 10693
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 5276 10733 5304 10764
rect 5534 10752 5540 10804
rect 5592 10752 5598 10804
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7469 10795 7527 10801
rect 7469 10792 7481 10795
rect 7156 10764 7481 10792
rect 7156 10752 7162 10764
rect 7469 10761 7481 10764
rect 7515 10792 7527 10795
rect 7650 10792 7656 10804
rect 7515 10764 7656 10792
rect 7515 10761 7527 10764
rect 7469 10755 7527 10761
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 9030 10752 9036 10804
rect 9088 10792 9094 10804
rect 9539 10795 9597 10801
rect 9539 10792 9551 10795
rect 9088 10764 9551 10792
rect 9088 10752 9094 10764
rect 9539 10761 9551 10764
rect 9585 10792 9597 10795
rect 15657 10795 15715 10801
rect 15657 10792 15669 10795
rect 9585 10764 9996 10792
rect 9585 10761 9597 10764
rect 9539 10755 9597 10761
rect 5261 10727 5319 10733
rect 5261 10693 5273 10727
rect 5307 10693 5319 10727
rect 9398 10724 9404 10736
rect 5261 10687 5319 10693
rect 7300 10696 7788 10724
rect 9154 10696 9404 10724
rect 2222 10616 2228 10668
rect 2280 10616 2286 10668
rect 4798 10616 4804 10668
rect 4856 10616 4862 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5031 10628 5457 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 5445 10625 5457 10628
rect 5491 10656 5503 10659
rect 5534 10656 5540 10668
rect 5491 10628 5540 10656
rect 5491 10625 5503 10628
rect 5445 10619 5503 10625
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10625 5871 10659
rect 5813 10619 5871 10625
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 6135 10628 6377 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 5721 10591 5779 10597
rect 5721 10588 5733 10591
rect 4948 10560 5733 10588
rect 4948 10548 4954 10560
rect 5721 10557 5733 10560
rect 5767 10557 5779 10591
rect 5721 10551 5779 10557
rect 5828 10520 5856 10619
rect 7006 10616 7012 10668
rect 7064 10616 7070 10668
rect 7300 10665 7328 10696
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10625 7159 10659
rect 7101 10619 7159 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6730 10588 6736 10600
rect 6227 10560 6736 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 7116 10588 7144 10619
rect 7466 10616 7472 10668
rect 7524 10616 7530 10668
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10656 7619 10659
rect 7760 10656 7788 10696
rect 9398 10684 9404 10696
rect 9456 10684 9462 10736
rect 8018 10656 8024 10668
rect 7607 10628 7696 10656
rect 7760 10628 8024 10656
rect 7607 10625 7619 10628
rect 7561 10619 7619 10625
rect 7484 10588 7512 10616
rect 7116 10560 7512 10588
rect 7558 10520 7564 10532
rect 5828 10492 7564 10520
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 5074 10412 5080 10464
rect 5132 10412 5138 10464
rect 7098 10412 7104 10464
rect 7156 10412 7162 10464
rect 7668 10452 7696 10628
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 9968 10665 9996 10764
rect 10704 10764 15669 10792
rect 10704 10668 10732 10764
rect 15657 10761 15669 10764
rect 15703 10761 15715 10795
rect 15657 10755 15715 10761
rect 16758 10752 16764 10804
rect 16816 10752 16822 10804
rect 19610 10792 19616 10804
rect 18800 10764 19616 10792
rect 10965 10727 11023 10733
rect 10965 10693 10977 10727
rect 11011 10724 11023 10727
rect 11330 10724 11336 10736
rect 11011 10696 11336 10724
rect 11011 10693 11023 10696
rect 10965 10687 11023 10693
rect 11330 10684 11336 10696
rect 11388 10724 11394 10736
rect 12618 10724 12624 10736
rect 11388 10696 12624 10724
rect 11388 10684 11394 10696
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 15194 10684 15200 10736
rect 15252 10684 15258 10736
rect 18800 10668 18828 10764
rect 19610 10752 19616 10764
rect 19668 10792 19674 10804
rect 19981 10795 20039 10801
rect 19981 10792 19993 10795
rect 19668 10764 19993 10792
rect 19668 10752 19674 10764
rect 19981 10761 19993 10764
rect 20027 10761 20039 10795
rect 19981 10755 20039 10761
rect 20165 10727 20223 10733
rect 20165 10724 20177 10727
rect 19720 10696 20177 10724
rect 19720 10668 19748 10696
rect 20165 10693 20177 10696
rect 20211 10693 20223 10727
rect 20165 10687 20223 10693
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 10192 10628 10425 10656
rect 10192 10616 10198 10628
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 10686 10616 10692 10668
rect 10744 10616 10750 10668
rect 10870 10616 10876 10668
rect 10928 10616 10934 10668
rect 11146 10665 11152 10668
rect 11109 10659 11152 10665
rect 11109 10625 11121 10659
rect 11109 10619 11152 10625
rect 11146 10616 11152 10619
rect 11204 10616 11210 10668
rect 11609 10659 11667 10665
rect 11609 10625 11621 10659
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10656 12127 10659
rect 12434 10656 12440 10668
rect 12115 10628 12440 10656
rect 12115 10625 12127 10628
rect 12069 10619 12127 10625
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 7926 10588 7932 10600
rect 7800 10560 7932 10588
rect 7800 10548 7806 10560
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8386 10588 8392 10600
rect 8159 10560 8392 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 11624 10588 11652 10619
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13872 10628 13921 10656
rect 13872 10616 13878 10628
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 17862 10616 17868 10668
rect 17920 10665 17926 10668
rect 17920 10656 17932 10665
rect 17920 10628 17965 10656
rect 17920 10619 17932 10628
rect 17920 10616 17926 10619
rect 18046 10616 18052 10668
rect 18104 10656 18110 10668
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 18104 10628 18153 10656
rect 18104 10616 18110 10628
rect 18141 10625 18153 10628
rect 18187 10656 18199 10659
rect 18233 10659 18291 10665
rect 18233 10656 18245 10659
rect 18187 10628 18245 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18233 10625 18245 10628
rect 18279 10625 18291 10659
rect 18233 10619 18291 10625
rect 18500 10659 18558 10665
rect 18500 10625 18512 10659
rect 18546 10656 18558 10659
rect 18782 10656 18788 10668
rect 18546 10628 18788 10656
rect 18546 10625 18558 10628
rect 18500 10619 18558 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 19702 10616 19708 10668
rect 19760 10616 19766 10668
rect 20070 10616 20076 10668
rect 20128 10616 20134 10668
rect 9876 10560 11652 10588
rect 9876 10532 9904 10560
rect 12158 10548 12164 10600
rect 12216 10548 12222 10600
rect 14182 10548 14188 10600
rect 14240 10548 14246 10600
rect 9858 10520 9864 10532
rect 9600 10492 9864 10520
rect 9600 10452 9628 10492
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 10229 10523 10287 10529
rect 10229 10520 10241 10523
rect 9968 10492 10241 10520
rect 9968 10464 9996 10492
rect 10229 10489 10241 10492
rect 10275 10489 10287 10523
rect 10229 10483 10287 10489
rect 11241 10523 11299 10529
rect 11241 10489 11253 10523
rect 11287 10520 11299 10523
rect 12176 10520 12204 10548
rect 19794 10520 19800 10532
rect 11287 10492 12204 10520
rect 19628 10492 19800 10520
rect 11287 10489 11299 10492
rect 11241 10483 11299 10489
rect 19628 10464 19656 10492
rect 19794 10480 19800 10492
rect 19852 10480 19858 10532
rect 7668 10424 9628 10452
rect 9674 10412 9680 10464
rect 9732 10412 9738 10464
rect 9950 10412 9956 10464
rect 10008 10412 10014 10464
rect 10042 10412 10048 10464
rect 10100 10412 10106 10464
rect 10137 10455 10195 10461
rect 10137 10421 10149 10455
rect 10183 10452 10195 10455
rect 10778 10452 10784 10464
rect 10183 10424 10784 10452
rect 10183 10421 10195 10424
rect 10137 10415 10195 10421
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11112 10424 11713 10452
rect 11112 10412 11118 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 13357 10455 13415 10461
rect 13357 10452 13369 10455
rect 13136 10424 13369 10452
rect 13136 10412 13142 10424
rect 13357 10421 13369 10424
rect 13403 10421 13415 10455
rect 13357 10415 13415 10421
rect 19610 10412 19616 10464
rect 19668 10412 19674 10464
rect 20349 10455 20407 10461
rect 20349 10421 20361 10455
rect 20395 10452 20407 10455
rect 20395 10424 20852 10452
rect 20395 10421 20407 10424
rect 20349 10415 20407 10421
rect 1104 10362 20792 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 10214 10362
rect 10266 10310 10278 10362
rect 10330 10310 10342 10362
rect 10394 10310 10406 10362
rect 10458 10310 10470 10362
rect 10522 10310 16214 10362
rect 16266 10310 16278 10362
rect 16330 10310 16342 10362
rect 16394 10310 16406 10362
rect 16458 10310 16470 10362
rect 16522 10310 20792 10362
rect 1104 10288 20792 10310
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 4798 10248 4804 10260
rect 3651 10220 4804 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 6641 10251 6699 10257
rect 6641 10217 6653 10251
rect 6687 10248 6699 10251
rect 7006 10248 7012 10260
rect 6687 10220 7012 10248
rect 6687 10217 6699 10220
rect 6641 10211 6699 10217
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 5552 10112 5580 10208
rect 6748 10121 6776 10220
rect 7006 10208 7012 10220
rect 7064 10248 7070 10260
rect 7742 10248 7748 10260
rect 7064 10220 7748 10248
rect 7064 10208 7070 10220
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 8481 10251 8539 10257
rect 8481 10248 8493 10251
rect 8076 10220 8493 10248
rect 8076 10208 8082 10220
rect 8481 10217 8493 10220
rect 8527 10217 8539 10251
rect 8481 10211 8539 10217
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8720 10220 8953 10248
rect 8720 10208 8726 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 9674 10208 9680 10260
rect 9732 10208 9738 10260
rect 9766 10208 9772 10260
rect 9824 10248 9830 10260
rect 10042 10248 10048 10260
rect 9824 10220 10048 10248
rect 9824 10208 9830 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 10689 10251 10747 10257
rect 10689 10248 10701 10251
rect 10652 10220 10701 10248
rect 10652 10208 10658 10220
rect 10689 10217 10701 10220
rect 10735 10217 10747 10251
rect 10689 10211 10747 10217
rect 13173 10251 13231 10257
rect 13173 10217 13185 10251
rect 13219 10248 13231 10251
rect 14182 10248 14188 10260
rect 13219 10220 14188 10248
rect 13219 10217 13231 10220
rect 13173 10211 13231 10217
rect 14182 10208 14188 10220
rect 14240 10208 14246 10260
rect 15749 10251 15807 10257
rect 15749 10217 15761 10251
rect 15795 10248 15807 10251
rect 15930 10248 15936 10260
rect 15795 10220 15936 10248
rect 15795 10217 15807 10220
rect 15749 10211 15807 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 18230 10208 18236 10260
rect 18288 10248 18294 10260
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 18288 10220 18429 10248
rect 18288 10208 18294 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 18417 10211 18475 10217
rect 20162 10208 20168 10260
rect 20220 10248 20226 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 20220 10220 20269 10248
rect 20220 10208 20226 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 1903 10084 3832 10112
rect 5552 10084 6193 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 3804 10053 3832 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10081 6791 10115
rect 6733 10075 6791 10081
rect 7466 10072 7472 10124
rect 7524 10112 7530 10124
rect 7742 10112 7748 10124
rect 7524 10084 7748 10112
rect 7524 10072 7530 10084
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 2133 9979 2191 9985
rect 2133 9945 2145 9979
rect 2179 9945 2191 9979
rect 3418 9976 3424 9988
rect 3358 9948 3424 9976
rect 2133 9939 2191 9945
rect 2148 9908 2176 9939
rect 3418 9936 3424 9948
rect 3476 9976 3482 9988
rect 3804 9976 3832 10007
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 9692 10044 9720 10208
rect 19610 10180 19616 10192
rect 18248 10152 19616 10180
rect 10870 10112 10876 10124
rect 10612 10084 10876 10112
rect 10612 10056 10640 10084
rect 10870 10072 10876 10084
rect 10928 10112 10934 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 10928 10084 11437 10112
rect 10928 10072 10934 10084
rect 11425 10081 11437 10084
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 9355 10016 9720 10044
rect 9769 10047 9827 10053
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 9769 10013 9781 10047
rect 9815 10044 9827 10047
rect 10505 10047 10563 10053
rect 10505 10044 10517 10047
rect 9815 10016 10517 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 10505 10013 10517 10016
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 3970 9976 3976 9988
rect 3476 9948 3740 9976
rect 3804 9948 3976 9976
rect 3476 9936 3482 9948
rect 2774 9908 2780 9920
rect 2148 9880 2780 9908
rect 2774 9868 2780 9880
rect 2832 9868 2838 9920
rect 3712 9908 3740 9948
rect 3970 9936 3976 9948
rect 4028 9936 4034 9988
rect 4065 9979 4123 9985
rect 4065 9945 4077 9979
rect 4111 9976 4123 9979
rect 4338 9976 4344 9988
rect 4111 9948 4344 9976
rect 4111 9945 4123 9948
rect 4065 9939 4123 9945
rect 4338 9936 4344 9948
rect 4396 9936 4402 9988
rect 4448 9948 4554 9976
rect 4448 9908 4476 9948
rect 6914 9936 6920 9988
rect 6972 9976 6978 9988
rect 7009 9979 7067 9985
rect 7009 9976 7021 9979
rect 6972 9948 7021 9976
rect 6972 9936 6978 9948
rect 7009 9945 7021 9948
rect 7055 9945 7067 9979
rect 7009 9939 7067 9945
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 9122 9976 9128 9988
rect 8812 9948 9128 9976
rect 8812 9936 8818 9948
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 3712 9880 4476 9908
rect 5626 9868 5632 9920
rect 5684 9868 5690 9920
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 8018 9908 8024 9920
rect 6696 9880 8024 9908
rect 6696 9868 6702 9880
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 9784 9908 9812 10007
rect 10594 10004 10600 10056
rect 10652 10004 10658 10056
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 11149 10047 11207 10053
rect 11149 10013 11161 10047
rect 11195 10013 11207 10047
rect 11149 10007 11207 10013
rect 9861 9979 9919 9985
rect 9861 9945 9873 9979
rect 9907 9976 9919 9979
rect 9950 9976 9956 9988
rect 9907 9948 9956 9976
rect 9907 9945 9919 9948
rect 9861 9939 9919 9945
rect 9950 9936 9956 9948
rect 10008 9976 10014 9988
rect 11164 9976 11192 10007
rect 11330 10004 11336 10056
rect 11388 10004 11394 10056
rect 13814 10004 13820 10056
rect 13872 10004 13878 10056
rect 14366 10004 14372 10056
rect 14424 10004 14430 10056
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 16761 10047 16819 10053
rect 16761 10044 16773 10047
rect 16172 10016 16773 10044
rect 16172 10004 16178 10016
rect 16761 10013 16773 10016
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 17028 10047 17086 10053
rect 17028 10013 17040 10047
rect 17074 10044 17086 10047
rect 18248 10044 18276 10152
rect 19610 10140 19616 10152
rect 19668 10140 19674 10192
rect 18877 10115 18935 10121
rect 18877 10081 18889 10115
rect 18923 10112 18935 10115
rect 20824 10112 20852 10424
rect 18923 10084 20852 10112
rect 18923 10081 18935 10084
rect 18877 10075 18935 10081
rect 17074 10016 18276 10044
rect 17074 10013 17086 10016
rect 17028 10007 17086 10013
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18601 10047 18659 10053
rect 18601 10044 18613 10047
rect 18380 10016 18613 10044
rect 18380 10004 18386 10016
rect 18601 10013 18613 10016
rect 18647 10013 18659 10047
rect 18601 10007 18659 10013
rect 18690 10004 18696 10056
rect 18748 10004 18754 10056
rect 19061 10047 19119 10053
rect 19061 10013 19073 10047
rect 19107 10044 19119 10047
rect 20162 10044 20168 10056
rect 19107 10016 20168 10044
rect 19107 10013 19119 10016
rect 19061 10007 19119 10013
rect 14642 9985 14648 9988
rect 10008 9948 11192 9976
rect 11241 9979 11299 9985
rect 10008 9936 10014 9948
rect 11241 9945 11253 9979
rect 11287 9976 11299 9979
rect 11701 9979 11759 9985
rect 11701 9976 11713 9979
rect 11287 9948 11713 9976
rect 11287 9945 11299 9948
rect 11241 9939 11299 9945
rect 11701 9945 11713 9948
rect 11747 9945 11759 9979
rect 13265 9979 13323 9985
rect 13265 9976 13277 9979
rect 12926 9948 13277 9976
rect 11701 9939 11759 9945
rect 13265 9945 13277 9948
rect 13311 9945 13323 9979
rect 14636 9976 14648 9985
rect 14603 9948 14648 9976
rect 13265 9939 13323 9945
rect 14636 9939 14648 9948
rect 14642 9936 14648 9939
rect 14700 9936 14706 9988
rect 18969 9979 19027 9985
rect 18969 9976 18981 9979
rect 18156 9948 18981 9976
rect 18156 9920 18184 9948
rect 18969 9945 18981 9948
rect 19015 9945 19027 9979
rect 18969 9939 19027 9945
rect 10042 9908 10048 9920
rect 9784 9880 10048 9908
rect 10042 9868 10048 9880
rect 10100 9868 10106 9920
rect 18138 9868 18144 9920
rect 18196 9868 18202 9920
rect 18230 9868 18236 9920
rect 18288 9908 18294 9920
rect 19076 9908 19104 10007
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 20349 10047 20407 10053
rect 20349 10013 20361 10047
rect 20395 10044 20407 10047
rect 20806 10044 20812 10056
rect 20395 10016 20812 10044
rect 20395 10013 20407 10016
rect 20349 10007 20407 10013
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 18288 9880 19104 9908
rect 18288 9868 18294 9880
rect 1104 9818 20792 9840
rect 1104 9766 7214 9818
rect 7266 9766 7278 9818
rect 7330 9766 7342 9818
rect 7394 9766 7406 9818
rect 7458 9766 7470 9818
rect 7522 9766 13214 9818
rect 13266 9766 13278 9818
rect 13330 9766 13342 9818
rect 13394 9766 13406 9818
rect 13458 9766 13470 9818
rect 13522 9766 19214 9818
rect 19266 9766 19278 9818
rect 19330 9766 19342 9818
rect 19394 9766 19406 9818
rect 19458 9766 19470 9818
rect 19522 9766 20792 9818
rect 1104 9744 20792 9766
rect 2774 9664 2780 9716
rect 2832 9664 2838 9716
rect 4338 9664 4344 9716
rect 4396 9664 4402 9716
rect 4890 9664 4896 9716
rect 4948 9664 4954 9716
rect 5074 9664 5080 9716
rect 5132 9664 5138 9716
rect 5626 9664 5632 9716
rect 5684 9664 5690 9716
rect 6822 9704 6828 9716
rect 6472 9676 6828 9704
rect 4356 9636 4384 9664
rect 4617 9639 4675 9645
rect 4617 9636 4629 9639
rect 4356 9608 4629 9636
rect 4617 9605 4629 9608
rect 4663 9605 4675 9639
rect 4908 9636 4936 9664
rect 4617 9599 4675 9605
rect 4816 9608 4936 9636
rect 4985 9639 5043 9645
rect 1578 9528 1584 9580
rect 1636 9568 1642 9580
rect 4816 9577 4844 9608
rect 4985 9605 4997 9639
rect 5031 9636 5043 9639
rect 5092 9636 5120 9664
rect 5644 9636 5672 9664
rect 6472 9636 6500 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 7469 9707 7527 9713
rect 7469 9704 7481 9707
rect 7300 9676 7481 9704
rect 5031 9608 5120 9636
rect 5276 9608 5672 9636
rect 5920 9608 6500 9636
rect 6549 9639 6607 9645
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 1765 9571 1823 9577
rect 1765 9568 1777 9571
rect 1636 9540 1777 9568
rect 1636 9528 1642 9540
rect 1765 9537 1777 9540
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 4157 9571 4215 9577
rect 3007 9540 3832 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3804 9441 3832 9540
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4801 9571 4859 9577
rect 4203 9540 4752 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9469 4491 9503
rect 4724 9500 4752 9540
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 4890 9528 4896 9580
rect 4948 9528 4954 9580
rect 4908 9500 4936 9528
rect 4724 9472 4936 9500
rect 5000 9500 5028 9599
rect 5074 9528 5080 9580
rect 5132 9577 5138 9580
rect 5276 9577 5304 9608
rect 5920 9580 5948 9608
rect 6549 9605 6561 9639
rect 6595 9636 6607 9639
rect 7098 9636 7104 9648
rect 6595 9608 7104 9636
rect 6595 9605 6607 9608
rect 6549 9599 6607 9605
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 5132 9571 5161 9577
rect 5149 9537 5161 9571
rect 5132 9531 5161 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 5132 9528 5138 9531
rect 5644 9500 5672 9531
rect 5902 9528 5908 9580
rect 5960 9528 5966 9580
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 5000 9472 5672 9500
rect 4433 9463 4491 9469
rect 3789 9435 3847 9441
rect 3789 9401 3801 9435
rect 3835 9401 3847 9435
rect 3789 9395 3847 9401
rect 1762 9324 1768 9376
rect 1820 9324 1826 9376
rect 3329 9367 3387 9373
rect 3329 9333 3341 9367
rect 3375 9364 3387 9367
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3375 9336 3709 9364
rect 3375 9333 3387 9336
rect 3329 9327 3387 9333
rect 3697 9333 3709 9336
rect 3743 9364 3755 9367
rect 3970 9364 3976 9376
rect 3743 9336 3976 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4264 9364 4292 9463
rect 4448 9432 4476 9463
rect 5718 9460 5724 9512
rect 5776 9460 5782 9512
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6380 9500 6408 9531
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7193 9571 7251 9577
rect 7193 9568 7205 9571
rect 7009 9531 7067 9537
rect 7116 9540 7205 9568
rect 7024 9500 7052 9531
rect 7116 9512 7144 9540
rect 7193 9537 7205 9540
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 5868 9472 7052 9500
rect 5868 9460 5874 9472
rect 7098 9460 7104 9512
rect 7156 9460 7162 9512
rect 4798 9432 4804 9444
rect 4448 9404 4804 9432
rect 4798 9392 4804 9404
rect 4856 9432 4862 9444
rect 5350 9432 5356 9444
rect 4856 9404 5356 9432
rect 4856 9392 4862 9404
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 6638 9432 6644 9444
rect 5920 9404 6644 9432
rect 4614 9364 4620 9376
rect 4264 9336 4620 9364
rect 4614 9324 4620 9336
rect 4672 9364 4678 9376
rect 5074 9364 5080 9376
rect 4672 9336 5080 9364
rect 4672 9324 4678 9336
rect 5074 9324 5080 9336
rect 5132 9364 5138 9376
rect 5442 9364 5448 9376
rect 5132 9336 5448 9364
rect 5132 9324 5138 9336
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5920 9373 5948 9404
rect 6638 9392 6644 9404
rect 6696 9392 6702 9444
rect 6730 9392 6736 9444
rect 6788 9432 6794 9444
rect 7300 9432 7328 9676
rect 7469 9673 7481 9676
rect 7515 9673 7527 9707
rect 7469 9667 7527 9673
rect 7558 9664 7564 9716
rect 7616 9664 7622 9716
rect 9766 9704 9772 9716
rect 9232 9676 9772 9704
rect 7377 9639 7435 9645
rect 7377 9605 7389 9639
rect 7423 9636 7435 9639
rect 7576 9636 7604 9664
rect 9232 9636 9260 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 10778 9704 10784 9716
rect 9916 9676 10784 9704
rect 9916 9664 9922 9676
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 12434 9664 12440 9716
rect 12492 9664 12498 9716
rect 18230 9704 18236 9716
rect 15120 9676 18236 9704
rect 14660 9648 14771 9674
rect 7423 9608 7604 9636
rect 7668 9608 9260 9636
rect 9335 9639 9393 9645
rect 7423 9605 7435 9608
rect 7377 9599 7435 9605
rect 7484 9509 7512 9608
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7668 9500 7696 9608
rect 9335 9605 9347 9639
rect 9381 9636 9393 9639
rect 9953 9639 10011 9645
rect 9953 9636 9965 9639
rect 9381 9608 9965 9636
rect 9381 9605 9393 9608
rect 9335 9599 9393 9605
rect 9953 9605 9965 9608
rect 9999 9605 10011 9639
rect 9953 9599 10011 9605
rect 14642 9596 14648 9648
rect 14700 9646 14771 9648
rect 14700 9596 14706 9646
rect 14743 9636 14771 9646
rect 15120 9636 15148 9676
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 18782 9664 18788 9716
rect 18840 9664 18846 9716
rect 14743 9608 15148 9636
rect 17420 9608 19012 9636
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 7926 9568 7932 9580
rect 7883 9540 7932 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 7469 9463 7527 9469
rect 7576 9472 7696 9500
rect 7760 9500 7788 9531
rect 7926 9528 7932 9540
rect 7984 9528 7990 9580
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 9030 9568 9036 9580
rect 8067 9540 9036 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8036 9500 8064 9531
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 7760 9472 8064 9500
rect 6788 9404 7328 9432
rect 6788 9392 6794 9404
rect 5905 9367 5963 9373
rect 5905 9364 5917 9367
rect 5684 9336 5917 9364
rect 5684 9324 5690 9336
rect 5905 9333 5917 9336
rect 5951 9333 5963 9367
rect 5905 9327 5963 9333
rect 6089 9367 6147 9373
rect 6089 9333 6101 9367
rect 6135 9364 6147 9367
rect 7576 9364 7604 9472
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8260 9472 8953 9500
rect 8260 9460 8266 9472
rect 8941 9469 8953 9472
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9232 9500 9260 9531
rect 9582 9528 9588 9580
rect 9640 9528 9646 9580
rect 10134 9528 10140 9580
rect 10192 9568 10198 9580
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 10192 9540 10517 9568
rect 10192 9528 10198 9540
rect 10505 9537 10517 9540
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 12345 9571 12403 9577
rect 12345 9537 12357 9571
rect 12391 9568 12403 9571
rect 12526 9568 12532 9580
rect 12391 9540 12532 9568
rect 12391 9537 12403 9540
rect 12345 9531 12403 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 14366 9528 14372 9580
rect 14424 9568 14430 9580
rect 14743 9577 14771 9608
rect 17420 9577 17448 9608
rect 14461 9571 14519 9577
rect 14461 9568 14473 9571
rect 14424 9540 14473 9568
rect 14424 9528 14430 9540
rect 14461 9537 14473 9540
rect 14507 9537 14519 9571
rect 14461 9531 14519 9537
rect 14728 9571 14786 9577
rect 14728 9537 14740 9571
rect 14774 9568 14786 9571
rect 17405 9571 17463 9577
rect 14774 9540 14808 9568
rect 14774 9537 14786 9540
rect 14728 9531 14786 9537
rect 17405 9537 17417 9571
rect 17451 9537 17463 9571
rect 17405 9531 17463 9537
rect 17672 9571 17730 9577
rect 17672 9537 17684 9571
rect 17718 9568 17730 9571
rect 17718 9540 18920 9568
rect 17718 9537 17730 9540
rect 17672 9531 17730 9537
rect 9232 9472 11284 9500
rect 7653 9435 7711 9441
rect 7653 9401 7665 9435
rect 7699 9432 7711 9435
rect 7926 9432 7932 9444
rect 7699 9404 7932 9432
rect 7699 9401 7711 9404
rect 7653 9395 7711 9401
rect 7926 9392 7932 9404
rect 7984 9432 7990 9444
rect 9030 9432 9036 9444
rect 7984 9404 9036 9432
rect 7984 9392 7990 9404
rect 9030 9392 9036 9404
rect 9088 9432 9094 9444
rect 9232 9432 9260 9472
rect 9088 9404 9260 9432
rect 9088 9392 9094 9404
rect 9306 9392 9312 9444
rect 9364 9432 9370 9444
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 9364 9404 9597 9432
rect 9364 9392 9370 9404
rect 9585 9401 9597 9404
rect 9631 9401 9643 9435
rect 9585 9395 9643 9401
rect 11256 9376 11284 9472
rect 6135 9336 7604 9364
rect 6135 9333 6147 9336
rect 6089 9327 6147 9333
rect 7834 9324 7840 9376
rect 7892 9324 7898 9376
rect 8389 9367 8447 9373
rect 8389 9333 8401 9367
rect 8435 9364 8447 9367
rect 8570 9364 8576 9376
rect 8435 9336 8576 9364
rect 8435 9333 8447 9336
rect 8389 9327 8447 9333
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 9272 9336 9505 9364
rect 9272 9324 9278 9336
rect 9493 9333 9505 9336
rect 9539 9333 9551 9367
rect 9493 9327 9551 9333
rect 11238 9324 11244 9376
rect 11296 9324 11302 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 12161 9367 12219 9373
rect 12161 9364 12173 9367
rect 11664 9336 12173 9364
rect 11664 9324 11670 9336
rect 12161 9333 12173 9336
rect 12207 9364 12219 9367
rect 15194 9364 15200 9376
rect 12207 9336 15200 9364
rect 12207 9333 12219 9336
rect 12161 9327 12219 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 15841 9367 15899 9373
rect 15841 9333 15853 9367
rect 15887 9364 15899 9367
rect 16574 9364 16580 9376
rect 15887 9336 16580 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 18892 9364 18920 9540
rect 18984 9512 19012 9608
rect 19236 9571 19294 9577
rect 19236 9537 19248 9571
rect 19282 9568 19294 9571
rect 19702 9568 19708 9580
rect 19282 9540 19708 9568
rect 19282 9537 19294 9540
rect 19236 9531 19294 9537
rect 19702 9528 19708 9540
rect 19760 9528 19766 9580
rect 18966 9460 18972 9512
rect 19024 9460 19030 9512
rect 20070 9364 20076 9376
rect 18892 9336 20076 9364
rect 20070 9324 20076 9336
rect 20128 9364 20134 9376
rect 20349 9367 20407 9373
rect 20349 9364 20361 9367
rect 20128 9336 20361 9364
rect 20128 9324 20134 9336
rect 20349 9333 20361 9336
rect 20395 9333 20407 9367
rect 20349 9327 20407 9333
rect 1104 9274 20792 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 10214 9274
rect 10266 9222 10278 9274
rect 10330 9222 10342 9274
rect 10394 9222 10406 9274
rect 10458 9222 10470 9274
rect 10522 9222 16214 9274
rect 16266 9222 16278 9274
rect 16330 9222 16342 9274
rect 16394 9222 16406 9274
rect 16458 9222 16470 9274
rect 16522 9222 20792 9274
rect 1104 9200 20792 9222
rect 1762 9120 1768 9172
rect 1820 9120 1826 9172
rect 5534 9120 5540 9172
rect 5592 9120 5598 9172
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 5810 9160 5816 9172
rect 5767 9132 5816 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 1780 8956 1808 9120
rect 5626 9024 5632 9036
rect 4816 8996 5632 9024
rect 4816 8965 4844 8996
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 1627 8928 1808 8956
rect 4801 8959 4859 8965
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 4801 8925 4813 8959
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5166 8956 5172 8968
rect 5123 8928 5172 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5166 8916 5172 8928
rect 5224 8956 5230 8968
rect 5736 8956 5764 9123
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 5902 9120 5908 9172
rect 5960 9120 5966 9172
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 7006 9160 7012 9172
rect 6963 9132 7012 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7742 9160 7748 9172
rect 7156 9132 7748 9160
rect 7156 9120 7162 9132
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 9122 9120 9128 9172
rect 9180 9120 9186 9172
rect 9214 9120 9220 9172
rect 9272 9120 9278 9172
rect 17770 9120 17776 9172
rect 17828 9120 17834 9172
rect 17865 9163 17923 9169
rect 17865 9129 17877 9163
rect 17911 9160 17923 9163
rect 18138 9160 18144 9172
rect 17911 9132 18144 9160
rect 17911 9129 17923 9132
rect 17865 9123 17923 9129
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 18233 9163 18291 9169
rect 18233 9129 18245 9163
rect 18279 9129 18291 9163
rect 18233 9123 18291 9129
rect 18417 9163 18475 9169
rect 18417 9129 18429 9163
rect 18463 9160 18475 9163
rect 18690 9160 18696 9172
rect 18463 9132 18696 9160
rect 18463 9129 18475 9132
rect 18417 9123 18475 9129
rect 5224 8928 5764 8956
rect 5224 8916 5230 8928
rect 4614 8848 4620 8900
rect 4672 8888 4678 8900
rect 4893 8891 4951 8897
rect 4893 8888 4905 8891
rect 4672 8860 4905 8888
rect 4672 8848 4678 8860
rect 4893 8857 4905 8860
rect 4939 8857 4951 8891
rect 4893 8851 4951 8857
rect 5350 8848 5356 8900
rect 5408 8848 5414 8900
rect 5569 8891 5627 8897
rect 5569 8857 5581 8891
rect 5615 8888 5627 8891
rect 5920 8888 5948 9120
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 7926 8956 7932 8968
rect 6328 8928 7932 8956
rect 6328 8916 6334 8928
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8260 8928 8953 8956
rect 8260 8916 8266 8928
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 9140 8956 9168 9120
rect 17589 9095 17647 9101
rect 17589 9061 17601 9095
rect 17635 9092 17647 9095
rect 18046 9092 18052 9104
rect 17635 9064 18052 9092
rect 17635 9061 17647 9064
rect 17589 9055 17647 9061
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 10134 9024 10140 9036
rect 9232 8996 10140 9024
rect 9232 8965 9260 8996
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 11054 9024 11060 9036
rect 10560 8996 11060 9024
rect 10560 8984 10566 8996
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 16574 9024 16580 9036
rect 12492 8996 13492 9024
rect 12492 8984 12498 8996
rect 8987 8928 9168 8956
rect 9217 8959 9275 8965
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9456 8928 9505 8956
rect 9456 8916 9462 8928
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 13464 8965 13492 8996
rect 16408 8996 16580 9024
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 11848 8928 13369 8956
rect 11848 8916 11854 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 16229 8959 16287 8965
rect 16229 8925 16241 8959
rect 16275 8956 16287 8959
rect 16408 8956 16436 8996
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 17957 9027 18015 9033
rect 17957 8993 17969 9027
rect 18003 9024 18015 9027
rect 18138 9024 18144 9036
rect 18003 8996 18144 9024
rect 18003 8993 18015 8996
rect 17957 8987 18015 8993
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 16275 8928 16436 8956
rect 16485 8959 16543 8965
rect 16275 8925 16287 8928
rect 16229 8919 16287 8925
rect 16485 8925 16497 8959
rect 16531 8956 16543 8959
rect 17678 8956 17684 8968
rect 16531 8928 17684 8956
rect 16531 8925 16543 8928
rect 16485 8919 16543 8925
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 18248 8956 18276 9123
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 17788 8928 18276 8956
rect 5615 8860 5948 8888
rect 5615 8857 5627 8860
rect 5569 8851 5627 8857
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 8297 8891 8355 8897
rect 8297 8888 8309 8891
rect 7616 8860 8309 8888
rect 7616 8848 7622 8860
rect 8297 8857 8309 8860
rect 8343 8857 8355 8891
rect 8297 8851 8355 8857
rect 8754 8848 8760 8900
rect 8812 8888 8818 8900
rect 8812 8860 9168 8888
rect 8812 8848 8818 8860
rect 2222 8780 2228 8832
rect 2280 8780 2286 8832
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4706 8820 4712 8832
rect 4304 8792 4712 8820
rect 4304 8780 4310 8792
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5258 8820 5264 8832
rect 5031 8792 5264 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 6454 8820 6460 8832
rect 5500 8792 6460 8820
rect 5500 8780 5506 8792
rect 6454 8780 6460 8792
rect 6512 8820 6518 8832
rect 7834 8820 7840 8832
rect 6512 8792 7840 8820
rect 6512 8780 6518 8792
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8076 8792 8401 8820
rect 8076 8780 8082 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 9030 8780 9036 8832
rect 9088 8780 9094 8832
rect 9140 8820 9168 8860
rect 9766 8848 9772 8900
rect 9824 8848 9830 8900
rect 10778 8848 10784 8900
rect 10836 8848 10842 8900
rect 11330 8848 11336 8900
rect 11388 8848 11394 8900
rect 12158 8848 12164 8900
rect 12216 8888 12222 8900
rect 13081 8891 13139 8897
rect 13081 8888 13093 8891
rect 12216 8860 13093 8888
rect 12216 8848 12222 8860
rect 13081 8857 13093 8860
rect 13127 8857 13139 8891
rect 13081 8851 13139 8857
rect 17586 8848 17592 8900
rect 17644 8848 17650 8900
rect 11146 8820 11152 8832
rect 9140 8792 11152 8820
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 11241 8823 11299 8829
rect 11241 8789 11253 8823
rect 11287 8820 11299 8823
rect 12066 8820 12072 8832
rect 11287 8792 12072 8820
rect 11287 8789 11299 8792
rect 11241 8783 11299 8789
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 13173 8823 13231 8829
rect 13173 8820 13185 8823
rect 12860 8792 13185 8820
rect 12860 8780 12866 8792
rect 13173 8789 13185 8792
rect 13219 8789 13231 8823
rect 13173 8783 13231 8789
rect 13538 8780 13544 8832
rect 13596 8780 13602 8832
rect 15105 8823 15163 8829
rect 15105 8789 15117 8823
rect 15151 8820 15163 8823
rect 15378 8820 15384 8832
rect 15151 8792 15384 8820
rect 15151 8789 15163 8792
rect 15105 8783 15163 8789
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 17788 8820 17816 8928
rect 18046 8848 18052 8900
rect 18104 8848 18110 8900
rect 17368 8792 17816 8820
rect 18259 8823 18317 8829
rect 17368 8780 17374 8792
rect 18259 8789 18271 8823
rect 18305 8820 18317 8823
rect 18782 8820 18788 8832
rect 18305 8792 18788 8820
rect 18305 8789 18317 8792
rect 18259 8783 18317 8789
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 1104 8730 20792 8752
rect 1104 8678 7214 8730
rect 7266 8678 7278 8730
rect 7330 8678 7342 8730
rect 7394 8678 7406 8730
rect 7458 8678 7470 8730
rect 7522 8678 13214 8730
rect 13266 8678 13278 8730
rect 13330 8678 13342 8730
rect 13394 8678 13406 8730
rect 13458 8678 13470 8730
rect 13522 8678 19214 8730
rect 19266 8678 19278 8730
rect 19330 8678 19342 8730
rect 19394 8678 19406 8730
rect 19458 8678 19470 8730
rect 19522 8678 20792 8730
rect 1104 8656 20792 8678
rect 2222 8576 2228 8628
rect 2280 8576 2286 8628
rect 5258 8616 5264 8628
rect 4172 8588 5264 8616
rect 2240 8480 2268 8576
rect 4172 8489 4200 8588
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5868 8588 5917 8616
rect 5868 8576 5874 8588
rect 5905 8585 5917 8588
rect 5951 8585 5963 8619
rect 5905 8579 5963 8585
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7064 8588 8033 8616
rect 7064 8576 7070 8588
rect 8021 8585 8033 8588
rect 8067 8616 8079 8619
rect 9306 8616 9312 8628
rect 8067 8588 8892 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 4246 8508 4252 8560
rect 4304 8508 4310 8560
rect 4430 8508 4436 8560
rect 4488 8557 4494 8560
rect 4488 8551 4517 8557
rect 4505 8517 4517 8551
rect 4488 8511 4517 8517
rect 4488 8508 4494 8511
rect 4706 8508 4712 8560
rect 4764 8508 4770 8560
rect 5721 8551 5779 8557
rect 5721 8548 5733 8551
rect 4908 8520 5733 8548
rect 4908 8489 4936 8520
rect 5721 8517 5733 8520
rect 5767 8548 5779 8551
rect 6733 8551 6791 8557
rect 5767 8520 5948 8548
rect 5767 8517 5779 8520
rect 5721 8511 5779 8517
rect 5920 8492 5948 8520
rect 6733 8517 6745 8551
rect 6779 8548 6791 8551
rect 6914 8548 6920 8560
rect 6779 8520 6920 8548
rect 6779 8517 6791 8520
rect 6733 8511 6791 8517
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7117 8551 7175 8557
rect 7117 8548 7129 8551
rect 7024 8520 7129 8548
rect 2409 8483 2467 8489
rect 2409 8480 2421 8483
rect 2240 8452 2421 8480
rect 2409 8449 2421 8452
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 4356 8412 4384 8443
rect 4356 8384 4476 8412
rect 4448 8344 4476 8384
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 4908 8412 4936 8443
rect 4672 8384 4936 8412
rect 4672 8372 4678 8384
rect 5092 8344 5120 8443
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 5537 8483 5595 8489
rect 5224 8452 5266 8480
rect 5224 8440 5230 8452
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 5626 8480 5632 8492
rect 5583 8452 5632 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6638 8480 6644 8492
rect 6595 8452 6644 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 6825 8483 6883 8489
rect 6825 8480 6837 8483
rect 6748 8452 6837 8480
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8412 6147 8415
rect 6748 8412 6776 8452
rect 6825 8449 6837 8452
rect 6871 8480 6883 8483
rect 7024 8480 7052 8520
rect 7117 8517 7129 8520
rect 7163 8517 7175 8551
rect 8202 8548 8208 8560
rect 7117 8511 7175 8517
rect 7576 8520 8208 8548
rect 7576 8489 7604 8520
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 8573 8551 8631 8557
rect 8573 8517 8585 8551
rect 8619 8548 8631 8551
rect 8754 8548 8760 8560
rect 8619 8520 8760 8548
rect 8619 8517 8631 8520
rect 8573 8511 8631 8517
rect 8754 8508 8760 8520
rect 8812 8508 8818 8560
rect 8864 8492 8892 8588
rect 9140 8588 9312 8616
rect 9140 8557 9168 8588
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 11258 8619 11316 8625
rect 9416 8588 10916 8616
rect 9416 8560 9444 8588
rect 9125 8551 9183 8557
rect 9125 8517 9137 8551
rect 9171 8517 9183 8551
rect 9125 8511 9183 8517
rect 9398 8508 9404 8560
rect 9456 8508 9462 8560
rect 10502 8548 10508 8560
rect 10350 8520 10508 8548
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 10888 8557 10916 8588
rect 11258 8585 11270 8619
rect 11304 8616 11316 8619
rect 12618 8616 12624 8628
rect 11304 8588 12624 8616
rect 11304 8585 11316 8588
rect 11258 8579 11316 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12802 8576 12808 8628
rect 12860 8576 12866 8628
rect 13538 8576 13544 8628
rect 13596 8616 13602 8628
rect 14001 8619 14059 8625
rect 13596 8588 13860 8616
rect 13596 8576 13602 8588
rect 10873 8551 10931 8557
rect 10873 8517 10885 8551
rect 10919 8517 10931 8551
rect 12434 8548 12440 8560
rect 10873 8511 10931 8517
rect 12268 8520 12440 8548
rect 6871 8452 7052 8480
rect 7561 8483 7619 8489
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 6135 8384 6776 8412
rect 6135 8381 6147 8384
rect 6089 8375 6147 8381
rect 6748 8356 6776 8384
rect 5626 8344 5632 8356
rect 4448 8316 4936 8344
rect 5092 8316 5632 8344
rect 4908 8288 4936 8316
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 6270 8304 6276 8356
rect 6328 8304 6334 8356
rect 6730 8304 6736 8356
rect 6788 8304 6794 8356
rect 7285 8347 7343 8353
rect 7285 8313 7297 8347
rect 7331 8344 7343 8347
rect 7576 8344 7604 8443
rect 8846 8440 8852 8492
rect 8904 8440 8910 8492
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 10962 8440 10968 8492
rect 11020 8440 11026 8492
rect 12268 8489 12296 8520
rect 12434 8508 12440 8520
rect 12492 8508 12498 8560
rect 12529 8551 12587 8557
rect 12529 8517 12541 8551
rect 12575 8548 12587 8551
rect 12820 8548 12848 8576
rect 12575 8520 12848 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 11085 8483 11143 8489
rect 11085 8449 11097 8483
rect 11131 8480 11143 8483
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 11131 8452 12265 8480
rect 11131 8449 11143 8452
rect 11085 8443 11143 8449
rect 12253 8449 12265 8452
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 13538 8440 13544 8492
rect 13596 8480 13602 8492
rect 13832 8480 13860 8588
rect 14001 8585 14013 8619
rect 14047 8585 14059 8619
rect 14001 8579 14059 8585
rect 14016 8548 14044 8579
rect 14274 8576 14280 8628
rect 14332 8616 14338 8628
rect 16393 8619 16451 8625
rect 14332 8588 14504 8616
rect 14332 8576 14338 8588
rect 14369 8551 14427 8557
rect 14369 8548 14381 8551
rect 14016 8520 14381 8548
rect 14369 8517 14381 8520
rect 14415 8517 14427 8551
rect 14476 8548 14504 8588
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 18046 8616 18052 8628
rect 16439 8588 18052 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18966 8576 18972 8628
rect 19024 8576 19030 8628
rect 19702 8576 19708 8628
rect 19760 8616 19766 8628
rect 19889 8619 19947 8625
rect 19889 8616 19901 8619
rect 19760 8588 19901 8616
rect 19760 8576 19766 8588
rect 19889 8585 19901 8588
rect 19935 8585 19947 8619
rect 19889 8579 19947 8585
rect 14476 8520 14858 8548
rect 14369 8511 14427 8517
rect 15930 8508 15936 8560
rect 15988 8548 15994 8560
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 15988 8520 16037 8548
rect 15988 8508 15994 8520
rect 16025 8517 16037 8520
rect 16071 8517 16083 8551
rect 16025 8511 16083 8517
rect 16241 8551 16299 8557
rect 16241 8517 16253 8551
rect 16287 8548 16299 8551
rect 16574 8548 16580 8560
rect 16287 8520 16580 8548
rect 16287 8517 16299 8520
rect 16241 8511 16299 8517
rect 16574 8508 16580 8520
rect 16632 8508 16638 8560
rect 18984 8548 19012 8576
rect 18524 8520 19012 8548
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13596 8452 13662 8480
rect 13832 8452 14105 8480
rect 13596 8440 13602 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 15896 8452 16681 8480
rect 15896 8440 15902 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 17678 8440 17684 8492
rect 17736 8480 17742 8492
rect 18524 8489 18552 8520
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 17736 8452 18429 8480
rect 17736 8440 17742 8452
rect 18417 8449 18429 8452
rect 18463 8480 18475 8483
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18463 8452 18521 8480
rect 18463 8449 18475 8452
rect 18417 8443 18475 8449
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18776 8483 18834 8489
rect 18776 8449 18788 8483
rect 18822 8480 18834 8483
rect 19058 8480 19064 8492
rect 18822 8452 19064 8480
rect 18822 8449 18834 8452
rect 18776 8443 18834 8449
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 11422 8412 11428 8424
rect 8772 8384 11428 8412
rect 8772 8353 8800 8384
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 11606 8372 11612 8424
rect 11664 8372 11670 8424
rect 12161 8415 12219 8421
rect 12161 8381 12173 8415
rect 12207 8381 12219 8415
rect 13814 8412 13820 8424
rect 12161 8375 12219 8381
rect 12360 8384 13820 8412
rect 7331 8316 7604 8344
rect 8205 8347 8263 8353
rect 7331 8313 7343 8316
rect 7285 8307 7343 8313
rect 8205 8313 8217 8347
rect 8251 8344 8263 8347
rect 8757 8347 8815 8353
rect 8251 8316 8708 8344
rect 8251 8313 8263 8316
rect 8205 8307 8263 8313
rect 1762 8236 1768 8288
rect 1820 8236 1826 8288
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3973 8279 4031 8285
rect 3973 8276 3985 8279
rect 3016 8248 3985 8276
rect 3016 8236 3022 8248
rect 3973 8245 3985 8248
rect 4019 8245 4031 8279
rect 3973 8239 4031 8245
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5166 8276 5172 8288
rect 4948 8248 5172 8276
rect 4948 8236 4954 8248
rect 5166 8236 5172 8248
rect 5224 8276 5230 8288
rect 6288 8276 6316 8304
rect 5224 8248 6316 8276
rect 5224 8236 5230 8248
rect 6362 8236 6368 8288
rect 6420 8236 6426 8288
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 7101 8279 7159 8285
rect 7101 8276 7113 8279
rect 6696 8248 7113 8276
rect 6696 8236 6702 8248
rect 7101 8245 7113 8248
rect 7147 8245 7159 8279
rect 7101 8239 7159 8245
rect 7466 8236 7472 8288
rect 7524 8236 7530 8288
rect 8386 8236 8392 8288
rect 8444 8276 8450 8288
rect 8573 8279 8631 8285
rect 8573 8276 8585 8279
rect 8444 8248 8585 8276
rect 8444 8236 8450 8248
rect 8573 8245 8585 8248
rect 8619 8245 8631 8279
rect 8680 8276 8708 8316
rect 8757 8313 8769 8347
rect 8803 8313 8815 8347
rect 8757 8307 8815 8313
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 10192 8316 10609 8344
rect 10192 8304 10198 8316
rect 10597 8313 10609 8316
rect 10643 8313 10655 8347
rect 12176 8344 12204 8375
rect 12360 8344 12388 8384
rect 13814 8372 13820 8384
rect 13872 8372 13878 8424
rect 12176 8316 12388 8344
rect 10597 8307 10655 8313
rect 15562 8304 15568 8356
rect 15620 8344 15626 8356
rect 15841 8347 15899 8353
rect 15841 8344 15853 8347
rect 15620 8316 15853 8344
rect 15620 8304 15626 8316
rect 15841 8313 15853 8316
rect 15887 8313 15899 8347
rect 15841 8307 15899 8313
rect 9858 8276 9864 8288
rect 8680 8248 9864 8276
rect 8573 8239 8631 8245
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 13078 8276 13084 8288
rect 12308 8248 13084 8276
rect 12308 8236 12314 8248
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 15378 8236 15384 8288
rect 15436 8276 15442 8288
rect 16022 8276 16028 8288
rect 15436 8248 16028 8276
rect 15436 8236 15442 8248
rect 16022 8236 16028 8248
rect 16080 8276 16086 8288
rect 16209 8279 16267 8285
rect 16209 8276 16221 8279
rect 16080 8248 16221 8276
rect 16080 8236 16086 8248
rect 16209 8245 16221 8248
rect 16255 8245 16267 8279
rect 16209 8239 16267 8245
rect 1104 8186 20792 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 10214 8186
rect 10266 8134 10278 8186
rect 10330 8134 10342 8186
rect 10394 8134 10406 8186
rect 10458 8134 10470 8186
rect 10522 8134 16214 8186
rect 16266 8134 16278 8186
rect 16330 8134 16342 8186
rect 16394 8134 16406 8186
rect 16458 8134 16470 8186
rect 16522 8134 20792 8186
rect 1104 8112 20792 8134
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 5537 8075 5595 8081
rect 3660 8044 5488 8072
rect 3660 8032 3666 8044
rect 5460 8004 5488 8044
rect 5537 8041 5549 8075
rect 5583 8072 5595 8075
rect 5810 8072 5816 8084
rect 5583 8044 5816 8072
rect 5583 8041 5595 8044
rect 5537 8035 5595 8041
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 9401 8075 9459 8081
rect 5920 8044 6592 8072
rect 5626 8004 5632 8016
rect 5460 7976 5632 8004
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 1762 7828 1768 7880
rect 1820 7828 1826 7880
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3651 7840 3801 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 5442 7868 5448 7880
rect 5198 7840 5448 7868
rect 3789 7831 3847 7837
rect 2498 7760 2504 7812
rect 2556 7760 2562 7812
rect 3804 7800 3832 7831
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 5920 7877 5948 8044
rect 6454 7964 6460 8016
rect 6512 7964 6518 8016
rect 6564 8004 6592 8044
rect 9401 8041 9413 8075
rect 9447 8072 9459 8075
rect 10594 8072 10600 8084
rect 9447 8044 10600 8072
rect 9447 8041 9459 8044
rect 9401 8035 9459 8041
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 10778 8032 10784 8084
rect 10836 8032 10842 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 10888 8044 13645 8072
rect 10888 8016 10916 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 16022 8032 16028 8084
rect 16080 8072 16086 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 16080 8044 16681 8072
rect 16080 8032 16086 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 17218 8032 17224 8084
rect 17276 8032 17282 8084
rect 17497 8075 17555 8081
rect 17497 8041 17509 8075
rect 17543 8072 17555 8075
rect 17586 8072 17592 8084
rect 17543 8044 17592 8072
rect 17543 8041 17555 8044
rect 17497 8035 17555 8041
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 18782 8032 18788 8084
rect 18840 8072 18846 8084
rect 19245 8075 19303 8081
rect 19245 8072 19257 8075
rect 18840 8044 19257 8072
rect 18840 8032 18846 8044
rect 19245 8041 19257 8044
rect 19291 8041 19303 8075
rect 19245 8035 19303 8041
rect 19352 8044 19932 8072
rect 7466 8004 7472 8016
rect 6564 7976 7472 8004
rect 7466 7964 7472 7976
rect 7524 7964 7530 8016
rect 10686 7964 10692 8016
rect 10744 8004 10750 8016
rect 10870 8004 10876 8016
rect 10744 7976 10876 8004
rect 10744 7964 10750 7976
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 11238 7964 11244 8016
rect 11296 8004 11302 8016
rect 11701 8007 11759 8013
rect 11701 8004 11713 8007
rect 11296 7976 11713 8004
rect 11296 7964 11302 7976
rect 11701 7973 11713 7976
rect 11747 7973 11759 8007
rect 11701 7967 11759 7973
rect 17037 8007 17095 8013
rect 17037 7973 17049 8007
rect 17083 8004 17095 8007
rect 18969 8007 19027 8013
rect 17083 7976 17264 8004
rect 17083 7973 17095 7976
rect 17037 7967 17095 7973
rect 6270 7936 6276 7948
rect 6104 7908 6276 7936
rect 6104 7877 6132 7908
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7936 6423 7939
rect 8757 7939 8815 7945
rect 6411 7908 6592 7936
rect 6411 7905 6423 7908
rect 6365 7899 6423 7905
rect 6564 7880 6592 7908
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 8846 7936 8852 7948
rect 8803 7908 8852 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 8846 7896 8852 7908
rect 8904 7896 8910 7948
rect 12250 7936 12256 7948
rect 10704 7908 12256 7936
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 6546 7828 6552 7880
rect 6604 7828 6610 7880
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7098 7868 7104 7880
rect 6963 7840 7104 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 10704 7877 10732 7908
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 17236 7945 17264 7976
rect 18969 7973 18981 8007
rect 19015 8004 19027 8007
rect 19058 8004 19064 8016
rect 19015 7976 19064 8004
rect 19015 7973 19027 7976
rect 18969 7967 19027 7973
rect 19058 7964 19064 7976
rect 19116 7964 19122 8016
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7905 17279 7939
rect 19352 7936 19380 8044
rect 19518 7964 19524 8016
rect 19576 8004 19582 8016
rect 19797 8007 19855 8013
rect 19797 8004 19809 8007
rect 19576 7976 19809 8004
rect 19576 7964 19582 7976
rect 19797 7973 19809 7976
rect 19843 7973 19855 8007
rect 19904 8004 19932 8044
rect 19978 8032 19984 8084
rect 20036 8032 20042 8084
rect 20349 8007 20407 8013
rect 20349 8004 20361 8007
rect 19904 7976 20361 8004
rect 19797 7967 19855 7973
rect 20349 7973 20361 7976
rect 20395 7973 20407 8007
rect 20349 7967 20407 7973
rect 17221 7899 17279 7905
rect 18708 7908 19380 7936
rect 19812 7936 19840 7967
rect 19812 7908 20208 7936
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 3970 7800 3976 7812
rect 3804 7772 3976 7800
rect 3970 7760 3976 7772
rect 4028 7760 4034 7812
rect 4062 7760 4068 7812
rect 4120 7760 4126 7812
rect 5350 7760 5356 7812
rect 5408 7800 5414 7812
rect 5721 7803 5779 7809
rect 5721 7800 5733 7803
rect 5408 7772 5733 7800
rect 5408 7760 5414 7772
rect 5721 7769 5733 7772
rect 5767 7769 5779 7803
rect 5721 7763 5779 7769
rect 5997 7803 6055 7809
rect 5997 7769 6009 7803
rect 6043 7769 6055 7803
rect 5997 7763 6055 7769
rect 6227 7803 6285 7809
rect 6227 7769 6239 7803
rect 6273 7800 6285 7803
rect 6472 7800 6500 7828
rect 6748 7800 6776 7828
rect 6273 7772 6500 7800
rect 6564 7772 6776 7800
rect 6273 7769 6285 7772
rect 6227 7763 6285 7769
rect 6012 7732 6040 7763
rect 6362 7732 6368 7744
rect 6012 7704 6368 7732
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 6454 7692 6460 7744
rect 6512 7732 6518 7744
rect 6564 7732 6592 7772
rect 8018 7760 8024 7812
rect 8076 7760 8082 7812
rect 8478 7760 8484 7812
rect 8536 7760 8542 7812
rect 10778 7760 10784 7812
rect 10836 7800 10842 7812
rect 11348 7800 11376 7831
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11480 7840 11529 7868
rect 11480 7828 11486 7840
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 15105 7871 15163 7877
rect 15105 7837 15117 7871
rect 15151 7868 15163 7871
rect 15194 7868 15200 7880
rect 15151 7840 15200 7868
rect 15151 7837 15163 7840
rect 15105 7831 15163 7837
rect 15194 7828 15200 7840
rect 15252 7868 15258 7880
rect 16114 7868 16120 7880
rect 15252 7840 16120 7868
rect 15252 7828 15258 7840
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16669 7871 16727 7877
rect 16669 7868 16681 7871
rect 16632 7840 16681 7868
rect 16632 7828 16638 7840
rect 16669 7837 16681 7840
rect 16715 7837 16727 7871
rect 16669 7831 16727 7837
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 17129 7871 17187 7877
rect 17129 7837 17141 7871
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 17678 7868 17684 7880
rect 17635 7840 17684 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 10836 7772 11560 7800
rect 10836 7760 10842 7772
rect 6512 7704 6592 7732
rect 6641 7735 6699 7741
rect 6512 7692 6518 7704
rect 6641 7701 6653 7735
rect 6687 7732 6699 7735
rect 6730 7732 6736 7744
rect 6687 7704 6736 7732
rect 6687 7701 6699 7704
rect 6641 7695 6699 7701
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 7006 7692 7012 7744
rect 7064 7692 7070 7744
rect 10686 7692 10692 7744
rect 10744 7732 10750 7744
rect 11422 7732 11428 7744
rect 10744 7704 11428 7732
rect 10744 7692 10750 7704
rect 11422 7692 11428 7704
rect 11480 7692 11486 7744
rect 11532 7732 11560 7772
rect 12066 7760 12072 7812
rect 12124 7800 12130 7812
rect 12161 7803 12219 7809
rect 12161 7800 12173 7803
rect 12124 7772 12173 7800
rect 12124 7760 12130 7772
rect 12161 7769 12173 7772
rect 12207 7769 12219 7803
rect 13538 7800 13544 7812
rect 13386 7772 13544 7800
rect 12161 7763 12219 7769
rect 13392 7732 13420 7772
rect 13538 7760 13544 7772
rect 13596 7800 13602 7812
rect 14274 7800 14280 7812
rect 13596 7772 14280 7800
rect 13596 7760 13602 7772
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 15378 7809 15384 7812
rect 15372 7800 15384 7809
rect 15339 7772 15384 7800
rect 15372 7763 15384 7772
rect 15378 7760 15384 7763
rect 15436 7760 15442 7812
rect 16776 7800 16804 7831
rect 16500 7772 16804 7800
rect 17144 7800 17172 7831
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 18708 7868 18736 7908
rect 17788 7840 18736 7868
rect 17788 7800 17816 7840
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 20180 7877 20208 7908
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 19116 7840 19533 7868
rect 19116 7828 19122 7840
rect 19521 7837 19533 7840
rect 19567 7868 19579 7871
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19567 7840 20085 7868
rect 19567 7837 19579 7840
rect 19521 7831 19579 7837
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 17144 7772 17816 7800
rect 17856 7803 17914 7809
rect 16500 7744 16528 7772
rect 17856 7769 17868 7803
rect 17902 7800 17914 7803
rect 18966 7800 18972 7812
rect 17902 7772 18972 7800
rect 17902 7769 17914 7772
rect 17856 7763 17914 7769
rect 18966 7760 18972 7772
rect 19024 7760 19030 7812
rect 19702 7800 19708 7812
rect 19536 7772 19708 7800
rect 11532 7704 13420 7732
rect 16482 7692 16488 7744
rect 16540 7692 16546 7744
rect 19429 7735 19487 7741
rect 19429 7701 19441 7735
rect 19475 7732 19487 7735
rect 19536 7732 19564 7772
rect 19702 7760 19708 7772
rect 19760 7800 19766 7812
rect 19889 7803 19947 7809
rect 19889 7800 19901 7803
rect 19760 7772 19901 7800
rect 19760 7760 19766 7772
rect 19889 7769 19901 7772
rect 19935 7769 19947 7803
rect 19889 7763 19947 7769
rect 19475 7704 19564 7732
rect 19613 7735 19671 7741
rect 19475 7701 19487 7704
rect 19429 7695 19487 7701
rect 19613 7701 19625 7735
rect 19659 7732 19671 7735
rect 19978 7732 19984 7744
rect 19659 7704 19984 7732
rect 19659 7701 19671 7704
rect 19613 7695 19671 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 1104 7642 20792 7664
rect 1104 7590 7214 7642
rect 7266 7590 7278 7642
rect 7330 7590 7342 7642
rect 7394 7590 7406 7642
rect 7458 7590 7470 7642
rect 7522 7590 13214 7642
rect 13266 7590 13278 7642
rect 13330 7590 13342 7642
rect 13394 7590 13406 7642
rect 13458 7590 13470 7642
rect 13522 7590 19214 7642
rect 19266 7590 19278 7642
rect 19330 7590 19342 7642
rect 19394 7590 19406 7642
rect 19458 7590 19470 7642
rect 19522 7590 20792 7642
rect 1104 7568 20792 7590
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4120 7500 4629 7528
rect 4120 7488 4126 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 5442 7528 5448 7540
rect 4617 7491 4675 7497
rect 4908 7500 5448 7528
rect 2685 7463 2743 7469
rect 2685 7429 2697 7463
rect 2731 7460 2743 7463
rect 2958 7460 2964 7472
rect 2731 7432 2964 7460
rect 2731 7429 2743 7432
rect 2685 7423 2743 7429
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 4908 7460 4936 7500
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 5626 7488 5632 7540
rect 5684 7488 5690 7540
rect 5718 7488 5724 7540
rect 5776 7488 5782 7540
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7528 6423 7531
rect 6546 7528 6552 7540
rect 6411 7500 6552 7528
rect 6411 7497 6423 7500
rect 6365 7491 6423 7497
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 7024 7500 8064 7528
rect 3910 7432 4936 7460
rect 4985 7463 5043 7469
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 5353 7463 5411 7469
rect 5353 7460 5365 7463
rect 5031 7432 5365 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 5353 7429 5365 7432
rect 5399 7429 5411 7463
rect 5644 7460 5672 7488
rect 7024 7460 7052 7500
rect 5644 7432 7052 7460
rect 5353 7423 5411 7429
rect 7098 7420 7104 7472
rect 7156 7460 7162 7472
rect 8036 7460 8064 7500
rect 8110 7488 8116 7540
rect 8168 7488 8174 7540
rect 8665 7531 8723 7537
rect 8665 7497 8677 7531
rect 8711 7528 8723 7531
rect 9398 7528 9404 7540
rect 8711 7500 9404 7528
rect 8711 7497 8723 7500
rect 8665 7491 8723 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 9508 7500 11468 7528
rect 7156 7432 7420 7460
rect 8036 7432 8340 7460
rect 7156 7420 7162 7432
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 4939 7364 5120 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 2409 7327 2467 7333
rect 2409 7324 2421 7327
rect 2332 7296 2421 7324
rect 2332 7200 2360 7296
rect 2409 7293 2421 7296
rect 2455 7293 2467 7327
rect 2409 7287 2467 7293
rect 4157 7327 4215 7333
rect 4157 7293 4169 7327
rect 4203 7324 4215 7327
rect 4614 7324 4620 7336
rect 4203 7296 4620 7324
rect 4203 7293 4215 7296
rect 4157 7287 4215 7293
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 4816 7324 4844 7355
rect 5092 7324 5120 7364
rect 5166 7352 5172 7404
rect 5224 7352 5230 7404
rect 5258 7352 5264 7404
rect 5316 7352 5322 7404
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5810 7392 5816 7404
rect 5491 7364 5816 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5460 7324 5488 7355
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6181 7395 6239 7401
rect 6181 7361 6193 7395
rect 6227 7392 6239 7395
rect 6270 7392 6276 7404
rect 6227 7364 6276 7392
rect 6227 7361 6239 7364
rect 6181 7355 6239 7361
rect 6270 7352 6276 7364
rect 6328 7392 6334 7404
rect 6638 7392 6644 7404
rect 6328 7364 6644 7392
rect 6328 7352 6334 7364
rect 6638 7352 6644 7364
rect 6696 7392 6702 7404
rect 7392 7401 7420 7432
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6696 7364 6929 7392
rect 6696 7352 6702 7364
rect 6917 7361 6929 7364
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 8312 7392 8340 7432
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 9508 7460 9536 7500
rect 8444 7432 9536 7460
rect 9953 7463 10011 7469
rect 8444 7420 8450 7432
rect 9953 7429 9965 7463
rect 9999 7460 10011 7463
rect 11330 7460 11336 7472
rect 9999 7432 11336 7460
rect 9999 7429 10011 7432
rect 9953 7423 10011 7429
rect 11330 7420 11336 7432
rect 11388 7420 11394 7472
rect 11440 7460 11468 7500
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 12437 7531 12495 7537
rect 12437 7528 12449 7531
rect 11940 7500 12449 7528
rect 11940 7488 11946 7500
rect 12437 7497 12449 7500
rect 12483 7497 12495 7531
rect 12437 7491 12495 7497
rect 17218 7488 17224 7540
rect 17276 7488 17282 7540
rect 18966 7488 18972 7540
rect 19024 7528 19030 7540
rect 19978 7528 19984 7540
rect 19024 7500 19984 7528
rect 19024 7488 19030 7500
rect 19978 7488 19984 7500
rect 20036 7488 20042 7540
rect 15930 7469 15936 7472
rect 15872 7463 15936 7469
rect 11440 7432 11928 7460
rect 7423 7364 8064 7392
rect 8312 7364 10640 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 4816 7296 4936 7324
rect 5092 7296 5488 7324
rect 4908 7256 4936 7296
rect 6086 7284 6092 7336
rect 6144 7324 6150 7336
rect 7006 7324 7012 7336
rect 6144 7296 7012 7324
rect 6144 7284 6150 7296
rect 7006 7284 7012 7296
rect 7064 7324 7070 7336
rect 7208 7324 7236 7355
rect 7064 7296 7236 7324
rect 7469 7327 7527 7333
rect 7064 7284 7070 7296
rect 7469 7293 7481 7327
rect 7515 7324 7527 7327
rect 7558 7324 7564 7336
rect 7515 7296 7564 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 6730 7256 6736 7268
rect 4908 7228 6736 7256
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 7098 7216 7104 7268
rect 7156 7256 7162 7268
rect 7484 7256 7512 7287
rect 7558 7284 7564 7296
rect 7616 7284 7622 7336
rect 7156 7228 7512 7256
rect 7156 7216 7162 7228
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 3970 7188 3976 7200
rect 2372 7160 3976 7188
rect 2372 7148 2378 7160
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5868 7160 5917 7188
rect 5868 7148 5874 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 5905 7151 5963 7157
rect 7374 7148 7380 7200
rect 7432 7148 7438 7200
rect 8036 7188 8064 7364
rect 10502 7216 10508 7268
rect 10560 7216 10566 7268
rect 10612 7256 10640 7364
rect 10686 7352 10692 7404
rect 10744 7352 10750 7404
rect 10870 7352 10876 7404
rect 10928 7352 10934 7404
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 11900 7401 11928 7432
rect 15872 7429 15884 7463
rect 15918 7429 15936 7463
rect 15872 7423 15936 7429
rect 15930 7420 15936 7423
rect 15988 7460 15994 7472
rect 16482 7460 16488 7472
rect 15988 7432 16488 7460
rect 15988 7420 15994 7432
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 18868 7463 18926 7469
rect 18868 7429 18880 7463
rect 18914 7460 18926 7463
rect 19058 7460 19064 7472
rect 18914 7432 19064 7460
rect 18914 7429 18926 7432
rect 18868 7423 18926 7429
rect 19058 7420 19064 7432
rect 19116 7420 19122 7472
rect 11609 7395 11667 7401
rect 11609 7392 11621 7395
rect 11020 7364 11621 7392
rect 11020 7352 11026 7364
rect 11609 7361 11621 7364
rect 11655 7361 11667 7395
rect 11609 7355 11667 7361
rect 11701 7395 11759 7401
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 12802 7392 12808 7404
rect 12575 7364 12808 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11716 7324 11744 7355
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 16114 7352 16120 7404
rect 16172 7352 16178 7404
rect 16761 7395 16819 7401
rect 16761 7392 16773 7395
rect 16224 7364 16773 7392
rect 11296 7296 11744 7324
rect 11296 7284 11302 7296
rect 10870 7256 10876 7268
rect 10612 7228 10876 7256
rect 10870 7216 10876 7228
rect 10928 7256 10934 7268
rect 11149 7259 11207 7265
rect 11149 7256 11161 7259
rect 10928 7228 11161 7256
rect 10928 7216 10934 7228
rect 11149 7225 11161 7228
rect 11195 7225 11207 7259
rect 11149 7219 11207 7225
rect 11333 7259 11391 7265
rect 11333 7225 11345 7259
rect 11379 7256 11391 7259
rect 11790 7256 11796 7268
rect 11379 7228 11796 7256
rect 11379 7225 11391 7228
rect 11333 7219 11391 7225
rect 11790 7216 11796 7228
rect 11848 7216 11854 7268
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 8036 7160 11713 7188
rect 11701 7157 11713 7160
rect 11747 7157 11759 7191
rect 11701 7151 11759 7157
rect 14737 7191 14795 7197
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 15470 7188 15476 7200
rect 14783 7160 15476 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 15470 7148 15476 7160
rect 15528 7188 15534 7200
rect 16224 7188 16252 7364
rect 16761 7361 16773 7364
rect 16807 7361 16819 7395
rect 16761 7355 16819 7361
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 17678 7352 17684 7404
rect 17736 7392 17742 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17736 7364 18613 7392
rect 17736 7352 17742 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 16853 7327 16911 7333
rect 16853 7324 16865 7327
rect 16632 7296 16865 7324
rect 16632 7284 16638 7296
rect 16853 7293 16865 7296
rect 16899 7293 16911 7327
rect 16853 7287 16911 7293
rect 15528 7160 16252 7188
rect 15528 7148 15534 7160
rect 16942 7148 16948 7200
rect 17000 7148 17006 7200
rect 1104 7098 20792 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 10214 7098
rect 10266 7046 10278 7098
rect 10330 7046 10342 7098
rect 10394 7046 10406 7098
rect 10458 7046 10470 7098
rect 10522 7046 16214 7098
rect 16266 7046 16278 7098
rect 16330 7046 16342 7098
rect 16394 7046 16406 7098
rect 16458 7046 16470 7098
rect 16522 7046 20792 7098
rect 1104 7024 20792 7046
rect 4788 6987 4846 6993
rect 4788 6953 4800 6987
rect 4834 6984 4846 6987
rect 5350 6984 5356 6996
rect 4834 6956 5356 6984
rect 4834 6953 4846 6956
rect 4788 6947 4846 6953
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 6270 6944 6276 6996
rect 6328 6944 6334 6996
rect 8386 6944 8392 6996
rect 8444 6944 8450 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10689 6987 10747 6993
rect 10689 6984 10701 6987
rect 9916 6956 10701 6984
rect 9916 6944 9922 6956
rect 10689 6953 10701 6956
rect 10735 6984 10747 6987
rect 10962 6984 10968 6996
rect 10735 6956 10968 6984
rect 10735 6953 10747 6956
rect 10689 6947 10747 6953
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 15194 6944 15200 6996
rect 15252 6944 15258 6996
rect 18969 6987 19027 6993
rect 18969 6953 18981 6987
rect 19015 6984 19027 6987
rect 19058 6984 19064 6996
rect 19015 6956 19064 6984
rect 19015 6953 19027 6956
rect 18969 6947 19027 6953
rect 19058 6944 19064 6956
rect 19116 6944 19122 6996
rect 8404 6916 8432 6944
rect 5920 6888 8064 6916
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 5920 6848 5948 6888
rect 8036 6860 8064 6888
rect 8312 6888 8432 6916
rect 5500 6820 5948 6848
rect 5500 6808 5506 6820
rect 3970 6740 3976 6792
rect 4028 6780 4034 6792
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4028 6752 4537 6780
rect 4028 6740 4034 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 5920 6766 5948 6820
rect 6564 6820 7420 6848
rect 4525 6743 4583 6749
rect 4433 6647 4491 6653
rect 4433 6613 4445 6647
rect 4479 6644 4491 6647
rect 4540 6644 4568 6743
rect 6086 6740 6092 6792
rect 6144 6740 6150 6792
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6454 6780 6460 6792
rect 6411 6752 6460 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 6564 6789 6592 6820
rect 7392 6792 7420 6820
rect 8018 6808 8024 6860
rect 8076 6808 8082 6860
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 6730 6740 6736 6792
rect 6788 6740 6794 6792
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8312 6780 8340 6888
rect 8260 6752 8340 6780
rect 8404 6820 8892 6848
rect 8260 6740 8266 6752
rect 6104 6712 6132 6740
rect 8404 6724 8432 6820
rect 8864 6792 8892 6820
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 15212 6857 15240 6944
rect 16761 6919 16819 6925
rect 16761 6885 16773 6919
rect 16807 6916 16819 6919
rect 17034 6916 17040 6928
rect 16807 6888 17040 6916
rect 16807 6885 16819 6888
rect 16761 6879 16819 6885
rect 17034 6876 17040 6888
rect 17092 6876 17098 6928
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 9824 6820 11069 6848
rect 9824 6808 9830 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6817 15255 6851
rect 15197 6811 15255 6817
rect 17310 6808 17316 6860
rect 17368 6808 17374 6860
rect 8478 6740 8484 6792
rect 8536 6740 8542 6792
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8904 6752 8953 6780
rect 8904 6740 8910 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10928 6752 10977 6780
rect 10928 6740 10934 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11146 6740 11152 6792
rect 11204 6740 11210 6792
rect 15470 6789 15476 6792
rect 15464 6780 15476 6789
rect 15431 6752 15476 6780
rect 15464 6743 15476 6752
rect 15528 6780 15534 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 15528 6752 17141 6780
rect 15470 6740 15476 6743
rect 15528 6740 15534 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 17129 6743 17187 6749
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6780 17647 6783
rect 17678 6780 17684 6792
rect 17635 6752 17684 6780
rect 17635 6749 17647 6752
rect 17589 6743 17647 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 6641 6715 6699 6721
rect 6641 6712 6653 6715
rect 6104 6684 6653 6712
rect 6641 6681 6653 6684
rect 6687 6681 6699 6715
rect 7009 6715 7067 6721
rect 7009 6712 7021 6715
rect 6641 6675 6699 6681
rect 6748 6684 7021 6712
rect 6748 6656 6776 6684
rect 7009 6681 7021 6684
rect 7055 6681 7067 6715
rect 7009 6675 7067 6681
rect 8021 6715 8079 6721
rect 8021 6681 8033 6715
rect 8067 6712 8079 6715
rect 8386 6712 8392 6724
rect 8067 6684 8392 6712
rect 8067 6681 8079 6684
rect 8021 6675 8079 6681
rect 8386 6672 8392 6684
rect 8444 6672 8450 6724
rect 5534 6644 5540 6656
rect 4479 6616 5540 6644
rect 4479 6613 4491 6616
rect 4433 6607 4491 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 6730 6604 6736 6656
rect 6788 6604 6794 6656
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 8496 6644 8524 6740
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 9217 6715 9275 6721
rect 9217 6712 9229 6715
rect 8803 6684 9229 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 9217 6681 9229 6684
rect 9263 6681 9275 6715
rect 10778 6712 10784 6724
rect 10442 6684 10784 6712
rect 9217 6675 9275 6681
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 11164 6712 11192 6740
rect 15562 6712 15568 6724
rect 11164 6684 15568 6712
rect 15562 6672 15568 6684
rect 15620 6672 15626 6724
rect 17037 6715 17095 6721
rect 17037 6712 17049 6715
rect 16868 6684 17049 6712
rect 6963 6616 8524 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 16868 6644 16896 6684
rect 17037 6681 17049 6684
rect 17083 6681 17095 6715
rect 17037 6675 17095 6681
rect 17856 6715 17914 6721
rect 17856 6681 17868 6715
rect 17902 6712 17914 6715
rect 19610 6712 19616 6724
rect 17902 6684 19616 6712
rect 17902 6681 17914 6684
rect 17856 6675 17914 6681
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 16632 6616 16896 6644
rect 16632 6604 16638 6616
rect 16942 6604 16948 6656
rect 17000 6604 17006 6656
rect 1104 6554 20792 6576
rect 1104 6502 7214 6554
rect 7266 6502 7278 6554
rect 7330 6502 7342 6554
rect 7394 6502 7406 6554
rect 7458 6502 7470 6554
rect 7522 6502 13214 6554
rect 13266 6502 13278 6554
rect 13330 6502 13342 6554
rect 13394 6502 13406 6554
rect 13458 6502 13470 6554
rect 13522 6502 19214 6554
rect 19266 6502 19278 6554
rect 19330 6502 19342 6554
rect 19394 6502 19406 6554
rect 19458 6502 19470 6554
rect 19522 6502 20792 6554
rect 1104 6480 20792 6502
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 8386 6440 8392 6452
rect 6227 6412 8392 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 2406 6332 2412 6384
rect 2464 6332 2470 6384
rect 5442 6372 5448 6384
rect 4278 6344 5448 6372
rect 2682 6264 2688 6316
rect 2740 6264 2746 6316
rect 1486 6196 1492 6248
rect 1544 6236 1550 6248
rect 1581 6239 1639 6245
rect 1581 6236 1593 6239
rect 1544 6208 1593 6236
rect 1544 6196 1550 6208
rect 1581 6205 1593 6208
rect 1627 6205 1639 6239
rect 1581 6199 1639 6205
rect 2774 6196 2780 6248
rect 2832 6196 2838 6248
rect 3050 6196 3056 6248
rect 3108 6196 3114 6248
rect 4062 6196 4068 6248
rect 4120 6236 4126 6248
rect 4356 6236 4384 6344
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 6380 6313 6408 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 12529 6443 12587 6449
rect 12529 6409 12541 6443
rect 12575 6409 12587 6443
rect 12529 6403 12587 6409
rect 14476 6412 14872 6440
rect 6641 6375 6699 6381
rect 6641 6341 6653 6375
rect 6687 6372 6699 6375
rect 6730 6372 6736 6384
rect 6687 6344 6736 6372
rect 6687 6341 6699 6344
rect 6641 6335 6699 6341
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 8018 6372 8024 6384
rect 7866 6344 8024 6372
rect 8018 6332 8024 6344
rect 8076 6332 8082 6384
rect 8202 6332 8208 6384
rect 8260 6332 8266 6384
rect 12544 6372 12572 6403
rect 12897 6375 12955 6381
rect 12897 6372 12909 6375
rect 12544 6344 12909 6372
rect 12897 6341 12909 6344
rect 12943 6341 12955 6375
rect 12897 6335 12955 6341
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5592 6276 6377 6304
rect 5592 6264 5598 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 4120 6208 4384 6236
rect 8113 6239 8171 6245
rect 4120 6196 4126 6208
rect 8113 6205 8125 6239
rect 8159 6236 8171 6239
rect 8220 6236 8248 6332
rect 9766 6264 9772 6316
rect 9824 6304 9830 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9824 6276 9965 6304
rect 9824 6264 9830 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 10045 6307 10103 6313
rect 10045 6273 10057 6307
rect 10091 6273 10103 6307
rect 10045 6267 10103 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 10962 6304 10968 6316
rect 10827 6276 10968 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 8159 6208 8248 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 10060 6236 10088 6267
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 9548 6208 10088 6236
rect 9548 6196 9554 6208
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 10192 6140 10701 6168
rect 10192 6128 10198 6140
rect 10689 6137 10701 6140
rect 10735 6137 10747 6171
rect 10689 6131 10747 6137
rect 11532 6112 11560 6267
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 11937 6307 11995 6313
rect 11937 6273 11949 6307
rect 11983 6304 11995 6307
rect 11983 6276 12296 6304
rect 11983 6273 11995 6276
rect 11937 6267 11995 6273
rect 2498 6060 2504 6112
rect 2556 6060 2562 6112
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4614 6100 4620 6112
rect 4571 6072 4620 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 8662 6060 8668 6112
rect 8720 6060 8726 6112
rect 10229 6103 10287 6109
rect 10229 6069 10241 6103
rect 10275 6100 10287 6103
rect 10778 6100 10784 6112
rect 10275 6072 10784 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 11514 6060 11520 6112
rect 11572 6060 11578 6112
rect 11808 6100 11836 6267
rect 12158 6236 12164 6248
rect 12084 6208 12164 6236
rect 12084 6177 12112 6208
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 12268 6236 12296 6276
rect 12342 6264 12348 6316
rect 12400 6264 12406 6316
rect 14366 6304 14372 6316
rect 14030 6276 14372 6304
rect 14366 6264 14372 6276
rect 14424 6304 14430 6316
rect 14476 6304 14504 6412
rect 14844 6372 14872 6412
rect 17034 6400 17040 6452
rect 17092 6440 17098 6452
rect 18049 6443 18107 6449
rect 18049 6440 18061 6443
rect 17092 6412 18061 6440
rect 17092 6400 17098 6412
rect 18049 6409 18061 6412
rect 18095 6409 18107 6443
rect 18049 6403 18107 6409
rect 18064 6372 18092 6403
rect 19610 6400 19616 6452
rect 19668 6400 19674 6452
rect 18478 6375 18536 6381
rect 18478 6372 18490 6375
rect 14844 6344 15226 6372
rect 16684 6344 17724 6372
rect 18064 6344 18490 6372
rect 16684 6313 16712 6344
rect 17696 6316 17724 6344
rect 18478 6341 18490 6344
rect 18524 6341 18536 6375
rect 18478 6335 18536 6341
rect 16942 6313 16948 6316
rect 14424 6276 14504 6304
rect 16669 6307 16727 6313
rect 14424 6264 14430 6276
rect 16669 6273 16681 6307
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 16936 6267 16948 6313
rect 17000 6304 17006 6316
rect 17310 6304 17316 6316
rect 17000 6276 17316 6304
rect 16942 6264 16948 6267
rect 17000 6264 17006 6276
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17678 6264 17684 6316
rect 17736 6304 17742 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17736 6276 18245 6304
rect 17736 6264 17742 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 12526 6236 12532 6248
rect 12268 6208 12532 6236
rect 12526 6196 12532 6208
rect 12584 6236 12590 6248
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12584 6208 12633 6236
rect 12584 6196 12590 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 14458 6196 14464 6248
rect 14516 6196 14522 6248
rect 14737 6239 14795 6245
rect 14737 6236 14749 6239
rect 14568 6208 14749 6236
rect 12069 6171 12127 6177
rect 12069 6137 12081 6171
rect 12115 6137 12127 6171
rect 12069 6131 12127 6137
rect 14369 6171 14427 6177
rect 14369 6137 14381 6171
rect 14415 6168 14427 6171
rect 14568 6168 14596 6208
rect 14737 6205 14749 6208
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 14415 6140 14596 6168
rect 14415 6137 14427 6140
rect 14369 6131 14427 6137
rect 14182 6100 14188 6112
rect 11808 6072 14188 6100
rect 14182 6060 14188 6072
rect 14240 6100 14246 6112
rect 16209 6103 16267 6109
rect 16209 6100 16221 6103
rect 14240 6072 16221 6100
rect 14240 6060 14246 6072
rect 16209 6069 16221 6072
rect 16255 6069 16267 6103
rect 16209 6063 16267 6069
rect 1104 6010 20792 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 10214 6010
rect 10266 5958 10278 6010
rect 10330 5958 10342 6010
rect 10394 5958 10406 6010
rect 10458 5958 10470 6010
rect 10522 5958 16214 6010
rect 16266 5958 16278 6010
rect 16330 5958 16342 6010
rect 16394 5958 16406 6010
rect 16458 5958 16470 6010
rect 16522 5958 20792 6010
rect 1104 5936 20792 5958
rect 2038 5896 2044 5908
rect 1688 5868 2044 5896
rect 1688 5769 1716 5868
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 3050 5856 3056 5908
rect 3108 5896 3114 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 3108 5868 3433 5896
rect 3108 5856 3114 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 3421 5859 3479 5865
rect 5534 5856 5540 5908
rect 5592 5856 5598 5908
rect 7377 5899 7435 5905
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 7558 5896 7564 5908
rect 7423 5868 7564 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 9033 5899 9091 5905
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9398 5896 9404 5908
rect 9079 5868 9404 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2498 5760 2504 5772
rect 1995 5732 2504 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 5552 5760 5580 5856
rect 5629 5763 5687 5769
rect 5629 5760 5641 5763
rect 5552 5732 5641 5760
rect 5629 5729 5641 5732
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 3602 5692 3608 5704
rect 3082 5664 3608 5692
rect 3602 5652 3608 5664
rect 3660 5692 3666 5704
rect 4062 5692 4068 5704
rect 3660 5664 4068 5692
rect 3660 5652 3666 5664
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 8294 5692 8300 5704
rect 7515 5664 8300 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 8941 5695 8999 5701
rect 8941 5661 8953 5695
rect 8987 5692 8999 5695
rect 9122 5692 9128 5704
rect 8987 5664 9128 5692
rect 8987 5661 8999 5664
rect 8941 5655 8999 5661
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9232 5701 9260 5868
rect 9398 5856 9404 5868
rect 9456 5856 9462 5908
rect 10134 5896 10140 5908
rect 9600 5868 10140 5896
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 9600 5760 9628 5868
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 10778 5856 10784 5908
rect 10836 5856 10842 5908
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 13633 5899 13691 5905
rect 13633 5896 13645 5899
rect 12400 5868 13645 5896
rect 12400 5856 12406 5868
rect 13633 5865 13645 5868
rect 13679 5865 13691 5899
rect 13633 5859 13691 5865
rect 14182 5856 14188 5908
rect 14240 5856 14246 5908
rect 17310 5856 17316 5908
rect 17368 5856 17374 5908
rect 9539 5732 9628 5760
rect 10796 5760 10824 5856
rect 13538 5788 13544 5840
rect 13596 5788 13602 5840
rect 13725 5831 13783 5837
rect 13725 5797 13737 5831
rect 13771 5797 13783 5831
rect 13725 5791 13783 5797
rect 13740 5760 13768 5791
rect 10796 5732 11376 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 5902 5584 5908 5636
rect 5960 5584 5966 5636
rect 8018 5624 8024 5636
rect 7130 5596 8024 5624
rect 8018 5584 8024 5596
rect 8076 5584 8082 5636
rect 8772 5624 8800 5652
rect 9416 5624 9444 5655
rect 10870 5652 10876 5704
rect 10928 5652 10934 5704
rect 11348 5701 11376 5732
rect 11532 5732 13768 5760
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5661 11391 5695
rect 11333 5655 11391 5661
rect 8772 5596 9444 5624
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 9769 5627 9827 5633
rect 9769 5624 9781 5627
rect 9732 5596 9781 5624
rect 9732 5584 9738 5596
rect 9769 5593 9781 5596
rect 9815 5593 9827 5627
rect 9769 5587 9827 5593
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 7653 5559 7711 5565
rect 7653 5525 7665 5559
rect 7699 5556 7711 5559
rect 8386 5556 8392 5568
rect 7699 5528 8392 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 9306 5516 9312 5568
rect 9364 5516 9370 5568
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 10888 5556 10916 5652
rect 11532 5624 11560 5732
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13596 5664 13737 5692
rect 13596 5652 13602 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5692 13967 5695
rect 14200 5692 14228 5856
rect 14553 5831 14611 5837
rect 14553 5797 14565 5831
rect 14599 5828 14611 5831
rect 14599 5800 15148 5828
rect 14599 5797 14611 5800
rect 14553 5791 14611 5797
rect 15120 5772 15148 5800
rect 15102 5720 15108 5772
rect 15160 5760 15166 5772
rect 15933 5763 15991 5769
rect 15933 5760 15945 5763
rect 15160 5732 15945 5760
rect 15160 5720 15166 5732
rect 15933 5729 15945 5732
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 13955 5664 14228 5692
rect 13955 5661 13967 5664
rect 13909 5655 13967 5661
rect 15838 5652 15844 5704
rect 15896 5652 15902 5704
rect 16200 5695 16258 5701
rect 16200 5661 16212 5695
rect 16246 5692 16258 5695
rect 16574 5692 16580 5704
rect 16246 5664 16580 5692
rect 16246 5661 16258 5664
rect 16200 5655 16258 5661
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 13173 5627 13231 5633
rect 13173 5624 13185 5627
rect 11164 5596 11560 5624
rect 12406 5596 13185 5624
rect 11164 5568 11192 5596
rect 9456 5528 10916 5556
rect 9456 5516 9462 5528
rect 11146 5516 11152 5568
rect 11204 5516 11210 5568
rect 11241 5559 11299 5565
rect 11241 5525 11253 5559
rect 11287 5556 11299 5559
rect 11514 5556 11520 5568
rect 11287 5528 11520 5556
rect 11287 5525 11299 5528
rect 11241 5519 11299 5525
rect 11514 5516 11520 5528
rect 11572 5556 11578 5568
rect 12406 5556 12434 5596
rect 13173 5593 13185 5596
rect 13219 5593 13231 5627
rect 13173 5587 13231 5593
rect 11572 5528 12434 5556
rect 11572 5516 11578 5528
rect 12618 5516 12624 5568
rect 12676 5516 12682 5568
rect 1104 5466 20792 5488
rect 1104 5414 7214 5466
rect 7266 5414 7278 5466
rect 7330 5414 7342 5466
rect 7394 5414 7406 5466
rect 7458 5414 7470 5466
rect 7522 5414 13214 5466
rect 13266 5414 13278 5466
rect 13330 5414 13342 5466
rect 13394 5414 13406 5466
rect 13458 5414 13470 5466
rect 13522 5414 19214 5466
rect 19266 5414 19278 5466
rect 19330 5414 19342 5466
rect 19394 5414 19406 5466
rect 19458 5414 19470 5466
rect 19522 5414 20792 5466
rect 1104 5392 20792 5414
rect 2038 5312 2044 5364
rect 2096 5312 2102 5364
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 2682 5352 2688 5364
rect 2547 5324 2688 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 2832 5324 3157 5352
rect 2832 5312 2838 5324
rect 3145 5321 3157 5324
rect 3191 5321 3203 5355
rect 3145 5315 3203 5321
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 4798 5352 4804 5364
rect 4387 5324 4804 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 7098 5352 7104 5364
rect 6472 5324 7104 5352
rect 1394 5176 1400 5228
rect 1452 5216 1458 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 1452 5188 1501 5216
rect 1452 5176 1458 5188
rect 1489 5185 1501 5188
rect 1535 5185 1547 5219
rect 2056 5216 2084 5312
rect 2314 5244 2320 5296
rect 2372 5244 2378 5296
rect 4614 5284 4620 5296
rect 3252 5256 3464 5284
rect 3252 5225 3280 5256
rect 3237 5219 3295 5225
rect 3237 5216 3249 5219
rect 2056 5188 3249 5216
rect 1489 5179 1547 5185
rect 3237 5185 3249 5188
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3142 5148 3148 5160
rect 3007 5120 3148 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 1578 5040 1584 5092
rect 1636 5080 1642 5092
rect 2593 5083 2651 5089
rect 2593 5080 2605 5083
rect 1636 5052 2605 5080
rect 1636 5040 1642 5052
rect 2593 5049 2605 5052
rect 2639 5080 2651 5083
rect 3344 5080 3372 5179
rect 3436 5148 3464 5256
rect 3804 5256 4620 5284
rect 3804 5225 3832 5256
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 3789 5219 3847 5225
rect 3789 5216 3801 5219
rect 3559 5188 3801 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3789 5185 3801 5188
rect 3835 5185 3847 5219
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3789 5179 3847 5185
rect 3896 5188 3985 5216
rect 3694 5148 3700 5160
rect 3436 5120 3700 5148
rect 3694 5108 3700 5120
rect 3752 5148 3758 5160
rect 3896 5148 3924 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4062 5176 4068 5228
rect 4120 5176 4126 5228
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 6472 5216 6500 5324
rect 7098 5312 7104 5324
rect 7156 5312 7162 5364
rect 8662 5312 8668 5364
rect 8720 5312 8726 5364
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9674 5352 9680 5364
rect 9263 5324 9680 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 12802 5312 12808 5364
rect 12860 5312 12866 5364
rect 14277 5355 14335 5361
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 14366 5352 14372 5364
rect 14323 5324 14372 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 14458 5312 14464 5364
rect 14516 5352 14522 5364
rect 14553 5355 14611 5361
rect 14553 5352 14565 5355
rect 14516 5324 14565 5352
rect 14516 5312 14522 5324
rect 14553 5321 14565 5324
rect 14599 5321 14611 5355
rect 14553 5315 14611 5321
rect 7116 5284 7144 5312
rect 7116 5256 7222 5284
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 8680 5284 8708 5312
rect 8352 5256 8616 5284
rect 8680 5256 8897 5284
rect 8352 5244 8358 5256
rect 5842 5188 6500 5216
rect 4157 5179 4215 5185
rect 3752 5120 3924 5148
rect 3752 5108 3758 5120
rect 2639 5052 3372 5080
rect 2639 5049 2651 5052
rect 2593 5043 2651 5049
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 4062 5080 4068 5092
rect 3476 5052 4068 5080
rect 3476 5040 3482 5052
rect 4062 5040 4068 5052
rect 4120 5080 4126 5092
rect 4172 5080 4200 5179
rect 8202 5176 8208 5228
rect 8260 5216 8266 5228
rect 8481 5219 8539 5225
rect 8481 5216 8493 5219
rect 8260 5188 8493 5216
rect 8260 5176 8266 5188
rect 8481 5185 8493 5188
rect 8527 5185 8539 5219
rect 8588 5216 8616 5256
rect 8869 5228 8897 5256
rect 9306 5244 9312 5296
rect 9364 5244 9370 5296
rect 10689 5287 10747 5293
rect 10689 5253 10701 5287
rect 10735 5284 10747 5287
rect 11146 5284 11152 5296
rect 10735 5256 11152 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 11517 5287 11575 5293
rect 11517 5284 11529 5287
rect 11388 5256 11529 5284
rect 11388 5244 11394 5256
rect 11517 5253 11529 5256
rect 11563 5253 11575 5287
rect 11517 5247 11575 5253
rect 13906 5244 13912 5296
rect 13964 5284 13970 5296
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 13964 5256 14197 5284
rect 13964 5244 13970 5256
rect 14185 5253 14197 5256
rect 14231 5253 14243 5287
rect 14185 5247 14243 5253
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 8588 5188 8677 5216
rect 8481 5179 8539 5185
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 8754 5176 8760 5228
rect 8812 5176 8818 5228
rect 8846 5176 8852 5228
rect 8904 5225 8910 5228
rect 8904 5219 8935 5225
rect 8923 5185 8935 5219
rect 8904 5179 8935 5185
rect 8904 5176 8910 5179
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5117 4491 5151
rect 4433 5111 4491 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4755 5120 6408 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4120 5052 4200 5080
rect 4120 5040 4126 5052
rect 3326 4972 3332 5024
rect 3384 4972 3390 5024
rect 4448 5012 4476 5111
rect 6380 5080 6408 5120
rect 6454 5108 6460 5160
rect 6512 5108 6518 5160
rect 9324 5148 9352 5244
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 9456 5188 9614 5216
rect 9456 5176 9462 5188
rect 11238 5176 11244 5228
rect 11296 5176 11302 5228
rect 14461 5219 14519 5225
rect 14461 5185 14473 5219
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5216 20499 5219
rect 20806 5216 20812 5228
rect 20487 5188 20812 5216
rect 20487 5185 20499 5188
rect 20441 5179 20499 5185
rect 6564 5120 9352 5148
rect 10965 5151 11023 5157
rect 6564 5080 6592 5120
rect 10965 5117 10977 5151
rect 11011 5117 11023 5151
rect 10965 5111 11023 5117
rect 6380 5052 6592 5080
rect 9033 5083 9091 5089
rect 9033 5049 9045 5083
rect 9079 5080 9091 5083
rect 9079 5052 9720 5080
rect 9079 5049 9091 5052
rect 9033 5043 9091 5049
rect 4706 5012 4712 5024
rect 4448 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6714 5015 6772 5021
rect 6714 5012 6726 5015
rect 6227 4984 6726 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6714 4981 6726 4984
rect 6760 4981 6772 5015
rect 6714 4975 6772 4981
rect 8202 4972 8208 5024
rect 8260 4972 8266 5024
rect 9692 5012 9720 5052
rect 10980 5012 11008 5111
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 13909 5151 13967 5157
rect 13909 5148 13921 5151
rect 12584 5120 13921 5148
rect 12584 5108 12590 5120
rect 13909 5117 13921 5120
rect 13955 5148 13967 5151
rect 14476 5148 14504 5179
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 13955 5120 14504 5148
rect 13955 5117 13967 5120
rect 13909 5111 13967 5117
rect 13262 5040 13268 5092
rect 13320 5080 13326 5092
rect 13320 5052 20300 5080
rect 13320 5040 13326 5052
rect 9692 4984 11008 5012
rect 11054 4972 11060 5024
rect 11112 4972 11118 5024
rect 13354 4972 13360 5024
rect 13412 4972 13418 5024
rect 20272 5021 20300 5052
rect 20257 5015 20315 5021
rect 20257 4981 20269 5015
rect 20303 4981 20315 5015
rect 20257 4975 20315 4981
rect 1104 4922 20792 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 10214 4922
rect 10266 4870 10278 4922
rect 10330 4870 10342 4922
rect 10394 4870 10406 4922
rect 10458 4870 10470 4922
rect 10522 4870 16214 4922
rect 16266 4870 16278 4922
rect 16330 4870 16342 4922
rect 16394 4870 16406 4922
rect 16458 4870 16470 4922
rect 16522 4870 20792 4922
rect 1104 4848 20792 4870
rect 4617 4811 4675 4817
rect 4617 4777 4629 4811
rect 4663 4808 4675 4811
rect 4706 4808 4712 4820
rect 4663 4780 4712 4808
rect 4663 4777 4675 4780
rect 4617 4771 4675 4777
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 4798 4768 4804 4820
rect 4856 4768 4862 4820
rect 5353 4811 5411 4817
rect 5353 4777 5365 4811
rect 5399 4808 5411 4811
rect 5902 4808 5908 4820
rect 5399 4780 5908 4808
rect 5399 4777 5411 4780
rect 5353 4771 5411 4777
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 6365 4811 6423 4817
rect 6365 4777 6377 4811
rect 6411 4808 6423 4811
rect 6454 4808 6460 4820
rect 6411 4780 6460 4808
rect 6411 4777 6423 4780
rect 6365 4771 6423 4777
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 12161 4811 12219 4817
rect 12161 4808 12173 4811
rect 11756 4780 12173 4808
rect 11756 4768 11762 4780
rect 12161 4777 12173 4780
rect 12207 4777 12219 4811
rect 13262 4808 13268 4820
rect 12161 4771 12219 4777
rect 12406 4780 13268 4808
rect 4080 4644 4660 4672
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 4080 4613 4108 4644
rect 4632 4616 4660 4644
rect 4065 4607 4123 4613
rect 3752 4576 3924 4604
rect 3752 4564 3758 4576
rect 3786 4496 3792 4548
rect 3844 4496 3850 4548
rect 3896 4536 3924 4576
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4212 4576 4445 4604
rect 4212 4564 4218 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4614 4564 4620 4616
rect 4672 4564 4678 4616
rect 4816 4604 4844 4768
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4816 4576 5273 4604
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5920 4604 5948 4768
rect 9122 4700 9128 4752
rect 9180 4740 9186 4752
rect 12406 4740 12434 4780
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13354 4768 13360 4820
rect 13412 4768 13418 4820
rect 9180 4712 12434 4740
rect 9180 4700 9186 4712
rect 6273 4607 6331 4613
rect 6273 4604 6285 4607
rect 5920 4576 6285 4604
rect 5261 4567 5319 4573
rect 6273 4573 6285 4576
rect 6319 4604 6331 4607
rect 8294 4604 8300 4616
rect 6319 4576 8300 4604
rect 6319 4573 6331 4576
rect 6273 4567 6331 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 9033 4607 9091 4613
rect 9033 4604 9045 4607
rect 8444 4576 9045 4604
rect 8444 4564 8450 4576
rect 9033 4573 9045 4576
rect 9079 4573 9091 4607
rect 12618 4604 12624 4616
rect 9033 4567 9091 4573
rect 12406 4576 12624 4604
rect 4249 4539 4307 4545
rect 4249 4536 4261 4539
rect 3896 4508 4261 4536
rect 4249 4505 4261 4508
rect 4295 4505 4307 4539
rect 4249 4499 4307 4505
rect 4341 4539 4399 4545
rect 4341 4505 4353 4539
rect 4387 4505 4399 4539
rect 8312 4536 8340 4564
rect 8478 4536 8484 4548
rect 8312 4508 8484 4536
rect 4341 4499 4399 4505
rect 3804 4468 3832 4496
rect 4356 4468 4384 4499
rect 8478 4496 8484 4508
rect 8536 4536 8542 4548
rect 9214 4536 9220 4548
rect 8536 4508 9220 4536
rect 8536 4496 8542 4508
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 10870 4496 10876 4548
rect 10928 4536 10934 4548
rect 12406 4536 12434 4576
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 13372 4604 13400 4768
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 13372 4576 13553 4604
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 13633 4607 13691 4613
rect 13633 4573 13645 4607
rect 13679 4573 13691 4607
rect 13633 4567 13691 4573
rect 13648 4536 13676 4567
rect 13814 4564 13820 4616
rect 13872 4564 13878 4616
rect 10928 4508 12434 4536
rect 13556 4508 13676 4536
rect 10928 4496 10934 4508
rect 13556 4480 13584 4508
rect 3804 4440 4384 4468
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 8754 4468 8760 4480
rect 8444 4440 8760 4468
rect 8444 4428 8450 4440
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 9766 4428 9772 4480
rect 9824 4468 9830 4480
rect 10321 4471 10379 4477
rect 10321 4468 10333 4471
rect 9824 4440 10333 4468
rect 9824 4428 9830 4440
rect 10321 4437 10333 4440
rect 10367 4437 10379 4471
rect 10321 4431 10379 4437
rect 12894 4428 12900 4480
rect 12952 4468 12958 4480
rect 13449 4471 13507 4477
rect 13449 4468 13461 4471
rect 12952 4440 13461 4468
rect 12952 4428 12958 4440
rect 13449 4437 13461 4440
rect 13495 4437 13507 4471
rect 13449 4431 13507 4437
rect 13538 4428 13544 4480
rect 13596 4428 13602 4480
rect 13722 4428 13728 4480
rect 13780 4428 13786 4480
rect 1104 4378 20792 4400
rect 1104 4326 7214 4378
rect 7266 4326 7278 4378
rect 7330 4326 7342 4378
rect 7394 4326 7406 4378
rect 7458 4326 7470 4378
rect 7522 4326 13214 4378
rect 13266 4326 13278 4378
rect 13330 4326 13342 4378
rect 13394 4326 13406 4378
rect 13458 4326 13470 4378
rect 13522 4326 19214 4378
rect 19266 4326 19278 4378
rect 19330 4326 19342 4378
rect 19394 4326 19406 4378
rect 19458 4326 19470 4378
rect 19522 4326 20792 4378
rect 1104 4304 20792 4326
rect 9122 4264 9128 4276
rect 8312 4236 9128 4264
rect 8312 4196 8340 4236
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 12897 4267 12955 4273
rect 12897 4264 12909 4267
rect 12584 4236 12909 4264
rect 12584 4224 12590 4236
rect 12897 4233 12909 4236
rect 12943 4233 12955 4267
rect 13722 4264 13728 4276
rect 12897 4227 12955 4233
rect 13372 4236 13728 4264
rect 8573 4199 8631 4205
rect 8573 4196 8585 4199
rect 8128 4168 8340 4196
rect 8404 4168 8585 4196
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3804 4100 3985 4128
rect 3804 4004 3832 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8128 4128 8156 4168
rect 8404 4140 8432 4168
rect 8573 4165 8585 4168
rect 8619 4165 8631 4199
rect 11054 4196 11060 4208
rect 8573 4159 8631 4165
rect 8864 4168 9449 4196
rect 8864 4140 8892 4168
rect 8067 4100 8156 4128
rect 8205 4131 8263 4137
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 8294 4128 8300 4140
rect 8251 4100 8300 4128
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8478 4088 8484 4140
rect 8536 4088 8542 4140
rect 8670 4131 8728 4137
rect 8670 4128 8682 4131
rect 8588 4100 8682 4128
rect 3786 3952 3792 4004
rect 3844 3952 3850 4004
rect 7024 3964 8156 3992
rect 7024 3936 7052 3964
rect 4062 3884 4068 3936
rect 4120 3884 4126 3936
rect 7006 3884 7012 3936
rect 7064 3884 7070 3936
rect 8018 3884 8024 3936
rect 8076 3884 8082 3936
rect 8128 3924 8156 3964
rect 8588 3924 8616 4100
rect 8670 4097 8682 4100
rect 8716 4097 8728 4131
rect 8670 4091 8728 4097
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9033 4131 9091 4137
rect 9033 4097 9045 4131
rect 9079 4128 9091 4131
rect 9122 4128 9128 4140
rect 9079 4100 9128 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9214 4088 9220 4140
rect 9272 4088 9278 4140
rect 9421 4137 9449 4168
rect 10888 4168 11060 4196
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9406 4131 9464 4137
rect 9406 4097 9418 4131
rect 9452 4128 9464 4131
rect 9582 4128 9588 4140
rect 9452 4100 9588 4128
rect 9452 4097 9464 4100
rect 9406 4091 9464 4097
rect 9324 4060 9352 4091
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 10220 4131 10278 4137
rect 10220 4097 10232 4131
rect 10266 4128 10278 4131
rect 10888 4128 10916 4168
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 13372 4205 13400 4236
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 13357 4199 13415 4205
rect 13357 4165 13369 4199
rect 13403 4165 13415 4199
rect 13357 4159 13415 4165
rect 14366 4156 14372 4208
rect 14424 4156 14430 4208
rect 10266 4100 10916 4128
rect 10266 4097 10278 4100
rect 10220 4091 10278 4097
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 11020 4100 11529 4128
rect 11020 4088 11026 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 11784 4131 11842 4137
rect 11784 4097 11796 4131
rect 11830 4128 11842 4131
rect 12894 4128 12900 4140
rect 11830 4100 12900 4128
rect 11830 4097 11842 4100
rect 11784 4091 11842 4097
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 9953 4063 10011 4069
rect 9953 4060 9965 4063
rect 9232 4032 9352 4060
rect 9692 4032 9965 4060
rect 9232 4004 9260 4032
rect 9214 3952 9220 4004
rect 9272 3952 9278 4004
rect 9490 3952 9496 4004
rect 9548 3992 9554 4004
rect 9585 3995 9643 4001
rect 9585 3992 9597 3995
rect 9548 3964 9597 3992
rect 9548 3952 9554 3964
rect 9585 3961 9597 3964
rect 9631 3961 9643 3995
rect 9585 3955 9643 3961
rect 9692 3936 9720 4032
rect 9953 4029 9965 4032
rect 9999 4029 10011 4063
rect 9953 4023 10011 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 8128 3896 8616 3924
rect 8846 3884 8852 3936
rect 8904 3884 8910 3936
rect 9674 3884 9680 3936
rect 9732 3884 9738 3936
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 12802 3924 12808 3936
rect 11379 3896 12808 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 12802 3884 12808 3896
rect 12860 3924 12866 3936
rect 13096 3924 13124 4023
rect 12860 3896 13124 3924
rect 12860 3884 12866 3896
rect 14826 3884 14832 3936
rect 14884 3884 14890 3936
rect 1104 3834 20792 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 10214 3834
rect 10266 3782 10278 3834
rect 10330 3782 10342 3834
rect 10394 3782 10406 3834
rect 10458 3782 10470 3834
rect 10522 3782 16214 3834
rect 16266 3782 16278 3834
rect 16330 3782 16342 3834
rect 16394 3782 16406 3834
rect 16458 3782 16470 3834
rect 16522 3782 20792 3834
rect 1104 3760 20792 3782
rect 14 3680 20 3732
rect 72 3720 78 3732
rect 1394 3720 1400 3732
rect 72 3692 1400 3720
rect 72 3680 78 3692
rect 1394 3680 1400 3692
rect 1452 3680 1458 3732
rect 3970 3680 3976 3732
rect 4028 3680 4034 3732
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 4120 3692 5764 3720
rect 4120 3680 4126 3692
rect 5736 3593 5764 3692
rect 8846 3680 8852 3732
rect 8904 3680 8910 3732
rect 9674 3680 9680 3732
rect 9732 3680 9738 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 12529 3723 12587 3729
rect 12529 3720 12541 3723
rect 12492 3692 12541 3720
rect 12492 3680 12498 3692
rect 12529 3689 12541 3692
rect 12575 3689 12587 3723
rect 13814 3720 13820 3732
rect 12529 3683 12587 3689
rect 13096 3692 13820 3720
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3553 5779 3587
rect 5721 3547 5779 3553
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 8018 3584 8024 3596
rect 7331 3556 8024 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 8864 3584 8892 3680
rect 12728 3624 13032 3652
rect 10229 3587 10287 3593
rect 10229 3584 10241 3587
rect 8352 3556 8708 3584
rect 8864 3556 10241 3584
rect 8352 3544 8358 3556
rect 3602 3476 3608 3528
rect 3660 3516 3666 3528
rect 4338 3516 4344 3528
rect 3660 3488 4344 3516
rect 3660 3476 3666 3488
rect 4338 3476 4344 3488
rect 4396 3476 4402 3528
rect 7006 3476 7012 3528
rect 7064 3476 7070 3528
rect 8570 3516 8576 3528
rect 8418 3488 8576 3516
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 8680 3516 8708 3556
rect 10229 3553 10241 3556
rect 10275 3553 10287 3587
rect 10229 3547 10287 3553
rect 9122 3516 9128 3528
rect 8680 3488 9128 3516
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9582 3525 9588 3528
rect 9401 3519 9459 3525
rect 9401 3516 9413 3519
rect 9272 3488 9413 3516
rect 9272 3476 9278 3488
rect 9401 3485 9413 3488
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 9545 3519 9588 3525
rect 9545 3485 9557 3519
rect 9545 3479 9588 3485
rect 9582 3476 9588 3479
rect 9640 3476 9646 3528
rect 12728 3525 12756 3624
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9692 3488 9873 3516
rect 5442 3408 5448 3460
rect 5500 3408 5506 3460
rect 7024 3380 7052 3476
rect 8680 3420 9260 3448
rect 8680 3380 8708 3420
rect 7024 3352 8708 3380
rect 8757 3383 8815 3389
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 8938 3380 8944 3392
rect 8803 3352 8944 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9232 3380 9260 3420
rect 9306 3408 9312 3460
rect 9364 3408 9370 3460
rect 9692 3380 9720 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 12345 3519 12403 3525
rect 12345 3485 12357 3519
rect 12391 3516 12403 3519
rect 12713 3519 12771 3525
rect 12391 3488 12425 3516
rect 12391 3485 12403 3488
rect 12345 3479 12403 3485
rect 12713 3485 12725 3519
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 10496 3451 10554 3457
rect 10496 3417 10508 3451
rect 10542 3448 10554 3451
rect 11514 3448 11520 3460
rect 10542 3420 11520 3448
rect 10542 3417 10554 3420
rect 10496 3411 10554 3417
rect 11514 3408 11520 3420
rect 11572 3408 11578 3460
rect 12360 3448 12388 3479
rect 12802 3476 12808 3528
rect 12860 3476 12866 3528
rect 12526 3448 12532 3460
rect 11624 3420 12532 3448
rect 9232 3352 9720 3380
rect 9950 3340 9956 3392
rect 10008 3340 10014 3392
rect 11624 3389 11652 3420
rect 12526 3408 12532 3420
rect 12584 3448 12590 3460
rect 12897 3451 12955 3457
rect 12897 3448 12909 3451
rect 12584 3420 12909 3448
rect 12584 3408 12590 3420
rect 12897 3417 12909 3420
rect 12943 3417 12955 3451
rect 13004 3448 13032 3624
rect 13096 3525 13124 3692
rect 13814 3680 13820 3692
rect 13872 3720 13878 3732
rect 14734 3720 14740 3732
rect 13872 3692 14740 3720
rect 13872 3680 13878 3692
rect 14734 3680 14740 3692
rect 14792 3680 14798 3732
rect 13538 3612 13544 3664
rect 13596 3612 13602 3664
rect 13633 3587 13691 3593
rect 13633 3553 13645 3587
rect 13679 3553 13691 3587
rect 13633 3547 13691 3553
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3584 14427 3587
rect 14826 3584 14832 3596
rect 14415 3556 14832 3584
rect 14415 3553 14427 3556
rect 14369 3547 14427 3553
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3485 13139 3519
rect 13648 3516 13676 3547
rect 14826 3544 14832 3556
rect 14884 3544 14890 3596
rect 13909 3519 13967 3525
rect 13909 3516 13921 3519
rect 13648 3488 13921 3516
rect 13081 3479 13139 3485
rect 13909 3485 13921 3488
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 14090 3476 14096 3528
rect 14148 3476 14154 3528
rect 13173 3451 13231 3457
rect 13173 3448 13185 3451
rect 13004 3420 13185 3448
rect 12897 3411 12955 3417
rect 13173 3417 13185 3420
rect 13219 3448 13231 3451
rect 13219 3420 13952 3448
rect 13219 3417 13231 3420
rect 13173 3411 13231 3417
rect 11609 3383 11667 3389
rect 11609 3349 11621 3383
rect 11655 3349 11667 3383
rect 11609 3343 11667 3349
rect 11790 3340 11796 3392
rect 11848 3340 11854 3392
rect 13722 3340 13728 3392
rect 13780 3340 13786 3392
rect 13924 3380 13952 3420
rect 14366 3408 14372 3460
rect 14424 3448 14430 3460
rect 14826 3448 14832 3460
rect 14424 3420 14832 3448
rect 14424 3408 14430 3420
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 15841 3383 15899 3389
rect 15841 3380 15853 3383
rect 13924 3352 15853 3380
rect 15841 3349 15853 3352
rect 15887 3349 15899 3383
rect 15841 3343 15899 3349
rect 1104 3290 20792 3312
rect 1104 3238 7214 3290
rect 7266 3238 7278 3290
rect 7330 3238 7342 3290
rect 7394 3238 7406 3290
rect 7458 3238 7470 3290
rect 7522 3238 13214 3290
rect 13266 3238 13278 3290
rect 13330 3238 13342 3290
rect 13394 3238 13406 3290
rect 13458 3238 13470 3290
rect 13522 3238 19214 3290
rect 19266 3238 19278 3290
rect 19330 3238 19342 3290
rect 19394 3238 19406 3290
rect 19458 3238 19470 3290
rect 19522 3238 20792 3290
rect 1104 3216 20792 3238
rect 5077 3179 5135 3185
rect 5077 3145 5089 3179
rect 5123 3176 5135 3179
rect 5442 3176 5448 3188
rect 5123 3148 5448 3176
rect 5123 3145 5135 3148
rect 5077 3139 5135 3145
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 8386 3136 8392 3188
rect 8444 3176 8450 3188
rect 8481 3179 8539 3185
rect 8481 3176 8493 3179
rect 8444 3148 8493 3176
rect 8444 3136 8450 3148
rect 8481 3145 8493 3148
rect 8527 3176 8539 3179
rect 9214 3176 9220 3188
rect 8527 3148 9220 3176
rect 8527 3145 8539 3148
rect 8481 3139 8539 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9950 3136 9956 3188
rect 10008 3136 10014 3188
rect 11514 3136 11520 3188
rect 11572 3136 11578 3188
rect 12710 3136 12716 3188
rect 12768 3136 12774 3188
rect 13722 3176 13728 3188
rect 12820 3148 13728 3176
rect 3326 3068 3332 3120
rect 3384 3108 3390 3120
rect 3605 3111 3663 3117
rect 3605 3108 3617 3111
rect 3384 3080 3617 3108
rect 3384 3068 3390 3080
rect 3605 3077 3617 3080
rect 3651 3077 3663 3111
rect 3605 3071 3663 3077
rect 4338 3068 4344 3120
rect 4396 3068 4402 3120
rect 9398 3068 9404 3120
rect 9456 3068 9462 3120
rect 9968 3108 9996 3136
rect 12728 3108 12756 3136
rect 12820 3117 12848 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 14792 3148 16129 3176
rect 14792 3136 14798 3148
rect 16117 3145 16129 3148
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 9968 3080 10272 3108
rect 8938 3000 8944 3052
rect 8996 3000 9002 3052
rect 10244 3049 10272 3080
rect 12268 3080 12756 3108
rect 12805 3111 12863 3117
rect 12268 3052 12296 3080
rect 12805 3077 12817 3111
rect 12851 3077 12863 3111
rect 14274 3108 14280 3120
rect 14030 3080 14280 3108
rect 12805 3071 12863 3077
rect 14274 3068 14280 3080
rect 14332 3108 14338 3120
rect 14332 3080 15134 3108
rect 14332 3068 14338 3080
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 12250 3000 12256 3052
rect 12308 3000 12314 3052
rect 12434 3000 12440 3052
rect 12492 3000 12498 3052
rect 12526 3000 12532 3052
rect 12584 3000 12590 3052
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 8956 2972 8984 3000
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 8956 2944 9965 2972
rect 3329 2935 3387 2941
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 9953 2935 10011 2941
rect 3344 2836 3372 2935
rect 10410 2932 10416 2984
rect 10468 2932 10474 2984
rect 10689 2975 10747 2981
rect 10689 2941 10701 2975
rect 10735 2941 10747 2975
rect 10689 2935 10747 2941
rect 3786 2836 3792 2848
rect 3344 2808 3792 2836
rect 3786 2796 3792 2808
rect 3844 2836 3850 2848
rect 10704 2836 10732 2935
rect 12066 2932 12072 2984
rect 12124 2932 12130 2984
rect 14366 2932 14372 2984
rect 14424 2932 14430 2984
rect 14645 2975 14703 2981
rect 14645 2972 14657 2975
rect 14476 2944 14657 2972
rect 14277 2907 14335 2913
rect 14277 2873 14289 2907
rect 14323 2904 14335 2907
rect 14476 2904 14504 2944
rect 14645 2941 14657 2944
rect 14691 2941 14703 2975
rect 14645 2935 14703 2941
rect 14323 2876 14504 2904
rect 14323 2873 14335 2876
rect 14277 2867 14335 2873
rect 20622 2864 20628 2916
rect 20680 2864 20686 2916
rect 3844 2808 10732 2836
rect 3844 2796 3850 2808
rect 12342 2796 12348 2848
rect 12400 2796 12406 2848
rect 13538 2796 13544 2848
rect 13596 2836 13602 2848
rect 20640 2836 20668 2864
rect 13596 2808 20668 2836
rect 13596 2796 13602 2808
rect 1104 2746 20792 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 10214 2746
rect 10266 2694 10278 2746
rect 10330 2694 10342 2746
rect 10394 2694 10406 2746
rect 10458 2694 10470 2746
rect 10522 2694 16214 2746
rect 16266 2694 16278 2746
rect 16330 2694 16342 2746
rect 16394 2694 16406 2746
rect 16458 2694 16470 2746
rect 16522 2694 20792 2746
rect 1104 2672 20792 2694
rect 9401 2635 9459 2641
rect 9401 2601 9413 2635
rect 9447 2632 9459 2635
rect 10962 2632 10968 2644
rect 9447 2604 10968 2632
rect 9447 2601 9459 2604
rect 9401 2595 9459 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 11977 2635 12035 2641
rect 11977 2601 11989 2635
rect 12023 2632 12035 2635
rect 12066 2632 12072 2644
rect 12023 2604 12072 2632
rect 12023 2601 12035 2604
rect 11977 2595 12035 2601
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12526 2592 12532 2644
rect 12584 2592 12590 2644
rect 13265 2635 13323 2641
rect 13265 2601 13277 2635
rect 13311 2632 13323 2635
rect 14366 2632 14372 2644
rect 13311 2604 14372 2632
rect 13311 2601 13323 2604
rect 13265 2595 13323 2601
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 5445 2567 5503 2573
rect 5445 2533 5457 2567
rect 5491 2564 5503 2567
rect 10042 2564 10048 2576
rect 5491 2536 10048 2564
rect 5491 2533 5503 2536
rect 5445 2527 5503 2533
rect 10042 2524 10048 2536
rect 10100 2524 10106 2576
rect 7006 2456 7012 2508
rect 7064 2456 7070 2508
rect 10965 2499 11023 2505
rect 10965 2465 10977 2499
rect 11011 2496 11023 2499
rect 11256 2496 11284 2592
rect 11011 2468 11284 2496
rect 11333 2499 11391 2505
rect 11011 2465 11023 2468
rect 10965 2459 11023 2465
rect 11333 2465 11345 2499
rect 11379 2496 11391 2499
rect 11609 2499 11667 2505
rect 11609 2496 11621 2499
rect 11379 2468 11621 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 11609 2465 11621 2468
rect 11655 2496 11667 2499
rect 12342 2496 12348 2508
rect 11655 2468 12348 2496
rect 11655 2465 11667 2468
rect 11609 2459 11667 2465
rect 12342 2456 12348 2468
rect 12400 2456 12406 2508
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 9766 2428 9772 2440
rect 8803 2400 9772 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 10870 2428 10876 2440
rect 10735 2400 10876 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2428 11759 2431
rect 11790 2428 11796 2440
rect 11747 2400 11796 2428
rect 11747 2397 11759 2400
rect 11701 2391 11759 2397
rect 11164 2360 11192 2391
rect 11790 2388 11796 2400
rect 11848 2388 11854 2440
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 12308 2400 12388 2428
rect 12308 2388 12314 2400
rect 12360 2369 12388 2400
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 12544 2428 12572 2592
rect 13633 2567 13691 2573
rect 13633 2533 13645 2567
rect 13679 2564 13691 2567
rect 14090 2564 14096 2576
rect 13679 2536 14096 2564
rect 13679 2533 13691 2536
rect 13633 2527 13691 2533
rect 14090 2524 14096 2536
rect 14148 2524 14154 2576
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12544 2400 13185 2428
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 12161 2363 12219 2369
rect 12161 2360 12173 2363
rect 11164 2332 12173 2360
rect 12161 2329 12173 2332
rect 12207 2329 12219 2363
rect 12161 2323 12219 2329
rect 12345 2363 12403 2369
rect 12345 2329 12357 2363
rect 12391 2329 12403 2363
rect 12452 2360 12480 2388
rect 12529 2363 12587 2369
rect 12529 2360 12541 2363
rect 12452 2332 12541 2360
rect 12345 2323 12403 2329
rect 12529 2329 12541 2332
rect 12575 2329 12587 2363
rect 12529 2323 12587 2329
rect 12360 2292 12388 2323
rect 13556 2292 13584 2391
rect 15194 2388 15200 2440
rect 15252 2428 15258 2440
rect 15749 2431 15807 2437
rect 15749 2428 15761 2431
rect 15252 2400 15761 2428
rect 15252 2388 15258 2400
rect 15749 2397 15761 2400
rect 15795 2397 15807 2431
rect 15749 2391 15807 2397
rect 15562 2320 15568 2372
rect 15620 2320 15626 2372
rect 12360 2264 13584 2292
rect 1104 2202 20792 2224
rect 1104 2150 7214 2202
rect 7266 2150 7278 2202
rect 7330 2150 7342 2202
rect 7394 2150 7406 2202
rect 7458 2150 7470 2202
rect 7522 2150 13214 2202
rect 13266 2150 13278 2202
rect 13330 2150 13342 2202
rect 13394 2150 13406 2202
rect 13458 2150 13470 2202
rect 13522 2150 19214 2202
rect 19266 2150 19278 2202
rect 19330 2150 19342 2202
rect 19394 2150 19406 2202
rect 19458 2150 19470 2202
rect 19522 2150 20792 2202
rect 1104 2128 20792 2150
<< via1 >>
rect 7214 21734 7266 21786
rect 7278 21734 7330 21786
rect 7342 21734 7394 21786
rect 7406 21734 7458 21786
rect 7470 21734 7522 21786
rect 13214 21734 13266 21786
rect 13278 21734 13330 21786
rect 13342 21734 13394 21786
rect 13406 21734 13458 21786
rect 13470 21734 13522 21786
rect 19214 21734 19266 21786
rect 19278 21734 19330 21786
rect 19342 21734 19394 21786
rect 19406 21734 19458 21786
rect 19470 21734 19522 21786
rect 3240 21496 3292 21548
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 13820 21564 13872 21616
rect 6920 21496 6972 21505
rect 5724 21428 5776 21480
rect 11520 21496 11572 21548
rect 18696 21496 18748 21548
rect 20260 21539 20312 21548
rect 20260 21505 20269 21539
rect 20269 21505 20303 21539
rect 20303 21505 20312 21539
rect 20260 21496 20312 21505
rect 10048 21471 10100 21480
rect 10048 21437 10057 21471
rect 10057 21437 10091 21471
rect 10091 21437 10100 21471
rect 10048 21428 10100 21437
rect 10876 21471 10928 21480
rect 10876 21437 10885 21471
rect 10885 21437 10919 21471
rect 10919 21437 10928 21471
rect 10876 21428 10928 21437
rect 7288 21335 7340 21344
rect 7288 21301 7297 21335
rect 7297 21301 7331 21335
rect 7331 21301 7340 21335
rect 7288 21292 7340 21301
rect 7564 21292 7616 21344
rect 7656 21292 7708 21344
rect 14280 21335 14332 21344
rect 14280 21301 14289 21335
rect 14289 21301 14323 21335
rect 14323 21301 14332 21335
rect 14280 21292 14332 21301
rect 18236 21292 18288 21344
rect 20444 21292 20496 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 10214 21190 10266 21242
rect 10278 21190 10330 21242
rect 10342 21190 10394 21242
rect 10406 21190 10458 21242
rect 10470 21190 10522 21242
rect 16214 21190 16266 21242
rect 16278 21190 16330 21242
rect 16342 21190 16394 21242
rect 16406 21190 16458 21242
rect 16470 21190 16522 21242
rect 7656 21131 7708 21140
rect 7656 21097 7665 21131
rect 7665 21097 7699 21131
rect 7699 21097 7708 21131
rect 7656 21088 7708 21097
rect 8392 21088 8444 21140
rect 10048 21088 10100 21140
rect 6276 20995 6328 21004
rect 6276 20961 6285 20995
rect 6285 20961 6319 20995
rect 6319 20961 6328 20995
rect 6276 20952 6328 20961
rect 7288 20952 7340 21004
rect 7564 20952 7616 21004
rect 4528 20791 4580 20800
rect 4528 20757 4537 20791
rect 4537 20757 4571 20791
rect 4571 20757 4580 20791
rect 4528 20748 4580 20757
rect 9588 20927 9640 20936
rect 9588 20893 9597 20927
rect 9597 20893 9631 20927
rect 9631 20893 9640 20927
rect 9588 20884 9640 20893
rect 8484 20748 8536 20800
rect 9404 20791 9456 20800
rect 9404 20757 9413 20791
rect 9413 20757 9447 20791
rect 9447 20757 9456 20791
rect 9404 20748 9456 20757
rect 9680 20748 9732 20800
rect 10876 20884 10928 20936
rect 13820 20884 13872 20936
rect 16120 20884 16172 20936
rect 12440 20748 12492 20800
rect 14556 20816 14608 20868
rect 17132 20816 17184 20868
rect 14280 20748 14332 20800
rect 17040 20748 17092 20800
rect 17868 20791 17920 20800
rect 17868 20757 17877 20791
rect 17877 20757 17911 20791
rect 17911 20757 17920 20791
rect 17868 20748 17920 20757
rect 7214 20646 7266 20698
rect 7278 20646 7330 20698
rect 7342 20646 7394 20698
rect 7406 20646 7458 20698
rect 7470 20646 7522 20698
rect 13214 20646 13266 20698
rect 13278 20646 13330 20698
rect 13342 20646 13394 20698
rect 13406 20646 13458 20698
rect 13470 20646 13522 20698
rect 19214 20646 19266 20698
rect 19278 20646 19330 20698
rect 19342 20646 19394 20698
rect 19406 20646 19458 20698
rect 19470 20646 19522 20698
rect 8484 20587 8536 20596
rect 8484 20553 8493 20587
rect 8493 20553 8527 20587
rect 8527 20553 8536 20587
rect 8484 20544 8536 20553
rect 17868 20544 17920 20596
rect 8300 20476 8352 20528
rect 11520 20476 11572 20528
rect 4528 20451 4580 20460
rect 4528 20417 4537 20451
rect 4537 20417 4571 20451
rect 4571 20417 4580 20451
rect 4528 20408 4580 20417
rect 13452 20451 13504 20460
rect 13820 20476 13872 20528
rect 13452 20417 13470 20451
rect 13470 20417 13504 20451
rect 13452 20408 13504 20417
rect 16764 20408 16816 20460
rect 17316 20408 17368 20460
rect 6276 20340 6328 20392
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 8392 20340 8444 20392
rect 10048 20383 10100 20392
rect 10048 20349 10057 20383
rect 10057 20349 10091 20383
rect 10091 20349 10100 20383
rect 10048 20340 10100 20349
rect 7012 20204 7064 20256
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 9680 20204 9732 20256
rect 16120 20383 16172 20392
rect 16120 20349 16129 20383
rect 16129 20349 16163 20383
rect 16163 20349 16172 20383
rect 16120 20340 16172 20349
rect 12348 20247 12400 20256
rect 12348 20213 12357 20247
rect 12357 20213 12391 20247
rect 12391 20213 12400 20247
rect 12348 20204 12400 20213
rect 14740 20247 14792 20256
rect 14740 20213 14749 20247
rect 14749 20213 14783 20247
rect 14783 20213 14792 20247
rect 14740 20204 14792 20213
rect 15384 20204 15436 20256
rect 17132 20204 17184 20256
rect 17960 20204 18012 20256
rect 19800 20204 19852 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 10214 20102 10266 20154
rect 10278 20102 10330 20154
rect 10342 20102 10394 20154
rect 10406 20102 10458 20154
rect 10470 20102 10522 20154
rect 16214 20102 16266 20154
rect 16278 20102 16330 20154
rect 16342 20102 16394 20154
rect 16406 20102 16458 20154
rect 16470 20102 16522 20154
rect 3884 20000 3936 20052
rect 6276 20000 6328 20052
rect 8392 20043 8444 20052
rect 8392 20009 8401 20043
rect 8401 20009 8435 20043
rect 8435 20009 8444 20043
rect 8392 20000 8444 20009
rect 10048 20000 10100 20052
rect 13452 20000 13504 20052
rect 14740 20000 14792 20052
rect 6920 19796 6972 19848
rect 9404 19864 9456 19916
rect 8576 19796 8628 19848
rect 11520 19796 11572 19848
rect 12440 19839 12492 19848
rect 12440 19805 12474 19839
rect 12474 19805 12492 19839
rect 12440 19796 12492 19805
rect 13636 19796 13688 19848
rect 14188 19839 14240 19848
rect 14188 19805 14197 19839
rect 14197 19805 14231 19839
rect 14231 19805 14240 19839
rect 14188 19796 14240 19805
rect 15292 19796 15344 19848
rect 6368 19771 6420 19780
rect 6368 19737 6377 19771
rect 6377 19737 6411 19771
rect 6411 19737 6420 19771
rect 6368 19728 6420 19737
rect 3516 19660 3568 19712
rect 6092 19660 6144 19712
rect 6184 19703 6236 19712
rect 6184 19669 6193 19703
rect 6193 19669 6227 19703
rect 6227 19669 6236 19703
rect 6184 19660 6236 19669
rect 7564 19660 7616 19712
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 17316 19796 17368 19848
rect 17040 19728 17092 19780
rect 17960 19796 18012 19848
rect 19800 19728 19852 19780
rect 17132 19703 17184 19712
rect 17132 19669 17141 19703
rect 17141 19669 17175 19703
rect 17175 19669 17184 19703
rect 17132 19660 17184 19669
rect 17408 19660 17460 19712
rect 17500 19703 17552 19712
rect 17500 19669 17509 19703
rect 17509 19669 17543 19703
rect 17543 19669 17552 19703
rect 17500 19660 17552 19669
rect 17684 19703 17736 19712
rect 17684 19669 17693 19703
rect 17693 19669 17727 19703
rect 17727 19669 17736 19703
rect 17684 19660 17736 19669
rect 7214 19558 7266 19610
rect 7278 19558 7330 19610
rect 7342 19558 7394 19610
rect 7406 19558 7458 19610
rect 7470 19558 7522 19610
rect 13214 19558 13266 19610
rect 13278 19558 13330 19610
rect 13342 19558 13394 19610
rect 13406 19558 13458 19610
rect 13470 19558 13522 19610
rect 19214 19558 19266 19610
rect 19278 19558 19330 19610
rect 19342 19558 19394 19610
rect 19406 19558 19458 19610
rect 19470 19558 19522 19610
rect 2780 19320 2832 19372
rect 3516 19320 3568 19372
rect 6276 19456 6328 19508
rect 6368 19456 6420 19508
rect 8576 19456 8628 19508
rect 11520 19456 11572 19508
rect 13084 19456 13136 19508
rect 7564 19431 7616 19440
rect 7564 19397 7582 19431
rect 7582 19397 7616 19431
rect 7564 19388 7616 19397
rect 4988 19363 5040 19372
rect 4988 19329 5022 19363
rect 5022 19329 5040 19363
rect 4988 19320 5040 19329
rect 9128 19320 9180 19372
rect 12348 19388 12400 19440
rect 13636 19388 13688 19440
rect 14188 19456 14240 19508
rect 16948 19456 17000 19508
rect 9588 19320 9640 19372
rect 16580 19388 16632 19440
rect 18052 19320 18104 19372
rect 18788 19363 18840 19372
rect 18788 19329 18822 19363
rect 18822 19329 18840 19363
rect 18788 19320 18840 19329
rect 7840 19295 7892 19304
rect 7840 19261 7849 19295
rect 7849 19261 7883 19295
rect 7883 19261 7892 19295
rect 7840 19252 7892 19261
rect 9312 19252 9364 19304
rect 9680 19252 9732 19304
rect 6184 19184 6236 19236
rect 8760 19184 8812 19236
rect 9220 19184 9272 19236
rect 11152 19295 11204 19304
rect 11152 19261 11161 19295
rect 11161 19261 11195 19295
rect 11195 19261 11204 19295
rect 11152 19252 11204 19261
rect 16672 19252 16724 19304
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 10048 19116 10100 19168
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 16856 19116 16908 19168
rect 17960 19159 18012 19168
rect 17960 19125 17969 19159
rect 17969 19125 18003 19159
rect 18003 19125 18012 19159
rect 17960 19116 18012 19125
rect 19892 19159 19944 19168
rect 19892 19125 19901 19159
rect 19901 19125 19935 19159
rect 19935 19125 19944 19159
rect 19892 19116 19944 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 10214 19014 10266 19066
rect 10278 19014 10330 19066
rect 10342 19014 10394 19066
rect 10406 19014 10458 19066
rect 10470 19014 10522 19066
rect 16214 19014 16266 19066
rect 16278 19014 16330 19066
rect 16342 19014 16394 19066
rect 16406 19014 16458 19066
rect 16470 19014 16522 19066
rect 4988 18912 5040 18964
rect 6368 18912 6420 18964
rect 6920 18912 6972 18964
rect 8760 18955 8812 18964
rect 8760 18921 8769 18955
rect 8769 18921 8803 18955
rect 8803 18921 8812 18955
rect 8760 18912 8812 18921
rect 9128 18912 9180 18964
rect 9588 18912 9640 18964
rect 11152 18912 11204 18964
rect 16764 18912 16816 18964
rect 16856 18955 16908 18964
rect 16856 18921 16865 18955
rect 16865 18921 16899 18955
rect 16899 18921 16908 18955
rect 16856 18912 16908 18921
rect 17132 18955 17184 18964
rect 17132 18921 17141 18955
rect 17141 18921 17175 18955
rect 17175 18921 17184 18955
rect 17132 18912 17184 18921
rect 18788 18912 18840 18964
rect 9496 18844 9548 18896
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 2780 18751 2832 18760
rect 2780 18717 2789 18751
rect 2789 18717 2823 18751
rect 2823 18717 2832 18751
rect 2780 18708 2832 18717
rect 6184 18751 6236 18760
rect 6184 18717 6193 18751
rect 6193 18717 6227 18751
rect 6227 18717 6236 18751
rect 6184 18708 6236 18717
rect 7012 18819 7064 18828
rect 7012 18785 7021 18819
rect 7021 18785 7055 18819
rect 7055 18785 7064 18819
rect 7012 18776 7064 18785
rect 7840 18776 7892 18828
rect 8300 18708 8352 18760
rect 8852 18776 8904 18828
rect 9312 18708 9364 18760
rect 7564 18640 7616 18692
rect 8576 18640 8628 18692
rect 9128 18640 9180 18692
rect 9772 18683 9824 18692
rect 9772 18649 9781 18683
rect 9781 18649 9815 18683
rect 9815 18649 9824 18683
rect 9772 18640 9824 18649
rect 2044 18615 2096 18624
rect 2044 18581 2053 18615
rect 2053 18581 2087 18615
rect 2087 18581 2096 18615
rect 2044 18572 2096 18581
rect 9404 18572 9456 18624
rect 11520 18776 11572 18828
rect 12348 18708 12400 18760
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 12992 18615 13044 18624
rect 12992 18581 13001 18615
rect 13001 18581 13035 18615
rect 13035 18581 13044 18615
rect 12992 18572 13044 18581
rect 15476 18640 15528 18692
rect 17040 18751 17092 18760
rect 17040 18717 17049 18751
rect 17049 18717 17083 18751
rect 17083 18717 17092 18751
rect 17040 18708 17092 18717
rect 17224 18708 17276 18760
rect 17408 18708 17460 18760
rect 17684 18708 17736 18760
rect 19892 18844 19944 18896
rect 17960 18640 18012 18692
rect 19616 18708 19668 18760
rect 19984 18683 20036 18692
rect 19984 18649 19993 18683
rect 19993 18649 20027 18683
rect 20027 18649 20036 18683
rect 19984 18640 20036 18649
rect 16120 18572 16172 18624
rect 19708 18615 19760 18624
rect 19708 18581 19717 18615
rect 19717 18581 19751 18615
rect 19751 18581 19760 18615
rect 19708 18572 19760 18581
rect 19800 18572 19852 18624
rect 7214 18470 7266 18522
rect 7278 18470 7330 18522
rect 7342 18470 7394 18522
rect 7406 18470 7458 18522
rect 7470 18470 7522 18522
rect 13214 18470 13266 18522
rect 13278 18470 13330 18522
rect 13342 18470 13394 18522
rect 13406 18470 13458 18522
rect 13470 18470 13522 18522
rect 19214 18470 19266 18522
rect 19278 18470 19330 18522
rect 19342 18470 19394 18522
rect 19406 18470 19458 18522
rect 19470 18470 19522 18522
rect 2044 18368 2096 18420
rect 7012 18368 7064 18420
rect 7564 18368 7616 18420
rect 9036 18368 9088 18420
rect 9220 18411 9272 18420
rect 9220 18377 9229 18411
rect 9229 18377 9263 18411
rect 9263 18377 9272 18411
rect 9220 18368 9272 18377
rect 9404 18368 9456 18420
rect 9772 18411 9824 18420
rect 9772 18377 9781 18411
rect 9781 18377 9815 18411
rect 9815 18377 9824 18411
rect 9772 18368 9824 18377
rect 9128 18300 9180 18352
rect 12992 18300 13044 18352
rect 13452 18300 13504 18352
rect 14280 18343 14332 18352
rect 14280 18309 14314 18343
rect 14314 18309 14332 18343
rect 14280 18300 14332 18309
rect 16672 18411 16724 18420
rect 16672 18377 16681 18411
rect 16681 18377 16715 18411
rect 16715 18377 16724 18411
rect 16672 18368 16724 18377
rect 15844 18300 15896 18352
rect 9496 18232 9548 18284
rect 10048 18232 10100 18284
rect 13820 18232 13872 18284
rect 16764 18232 16816 18284
rect 19708 18368 19760 18420
rect 9588 18164 9640 18216
rect 19432 18300 19484 18352
rect 19892 18300 19944 18352
rect 9496 18096 9548 18148
rect 2136 18071 2188 18080
rect 2136 18037 2145 18071
rect 2145 18037 2179 18071
rect 2179 18037 2188 18071
rect 2136 18028 2188 18037
rect 9312 18028 9364 18080
rect 12532 18071 12584 18080
rect 12532 18037 12541 18071
rect 12541 18037 12575 18071
rect 12575 18037 12584 18071
rect 12532 18028 12584 18037
rect 13176 18028 13228 18080
rect 15476 18028 15528 18080
rect 17500 18028 17552 18080
rect 17592 18071 17644 18080
rect 17592 18037 17601 18071
rect 17601 18037 17635 18071
rect 17635 18037 17644 18071
rect 17592 18028 17644 18037
rect 17960 18096 18012 18148
rect 19708 18028 19760 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 10214 17926 10266 17978
rect 10278 17926 10330 17978
rect 10342 17926 10394 17978
rect 10406 17926 10458 17978
rect 10470 17926 10522 17978
rect 16214 17926 16266 17978
rect 16278 17926 16330 17978
rect 16342 17926 16394 17978
rect 16406 17926 16458 17978
rect 16470 17926 16522 17978
rect 12624 17824 12676 17876
rect 13452 17824 13504 17876
rect 15476 17824 15528 17876
rect 18052 17824 18104 17876
rect 19616 17867 19668 17876
rect 19616 17833 19625 17867
rect 19625 17833 19659 17867
rect 19659 17833 19668 17867
rect 19616 17824 19668 17833
rect 18604 17756 18656 17808
rect 1676 17620 1728 17672
rect 2688 17552 2740 17604
rect 1400 17484 1452 17536
rect 3792 17663 3844 17672
rect 3792 17629 3801 17663
rect 3801 17629 3835 17663
rect 3835 17629 3844 17663
rect 3792 17620 3844 17629
rect 4804 17620 4856 17672
rect 5356 17663 5408 17672
rect 5356 17629 5365 17663
rect 5365 17629 5399 17663
rect 5399 17629 5408 17663
rect 5356 17620 5408 17629
rect 6092 17688 6144 17740
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 17960 17688 18012 17740
rect 19984 17688 20036 17740
rect 11520 17620 11572 17672
rect 13728 17620 13780 17672
rect 15844 17663 15896 17672
rect 15844 17629 15862 17663
rect 15862 17629 15896 17663
rect 15844 17620 15896 17629
rect 16948 17620 17000 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 19800 17620 19852 17672
rect 12532 17552 12584 17604
rect 12900 17552 12952 17604
rect 13176 17552 13228 17604
rect 13452 17595 13504 17604
rect 13452 17561 13461 17595
rect 13461 17561 13495 17595
rect 13495 17561 13504 17595
rect 13452 17552 13504 17561
rect 14280 17552 14332 17604
rect 18052 17552 18104 17604
rect 4252 17484 4304 17536
rect 4620 17527 4672 17536
rect 4620 17493 4629 17527
rect 4629 17493 4663 17527
rect 4663 17493 4672 17527
rect 4620 17484 4672 17493
rect 5080 17484 5132 17536
rect 5540 17484 5592 17536
rect 5632 17527 5684 17536
rect 5632 17493 5641 17527
rect 5641 17493 5675 17527
rect 5675 17493 5684 17527
rect 5632 17484 5684 17493
rect 11428 17484 11480 17536
rect 11612 17527 11664 17536
rect 11612 17493 11621 17527
rect 11621 17493 11655 17527
rect 11655 17493 11664 17527
rect 11612 17484 11664 17493
rect 12992 17484 13044 17536
rect 13544 17484 13596 17536
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 7214 17382 7266 17434
rect 7278 17382 7330 17434
rect 7342 17382 7394 17434
rect 7406 17382 7458 17434
rect 7470 17382 7522 17434
rect 13214 17382 13266 17434
rect 13278 17382 13330 17434
rect 13342 17382 13394 17434
rect 13406 17382 13458 17434
rect 13470 17382 13522 17434
rect 19214 17382 19266 17434
rect 19278 17382 19330 17434
rect 19342 17382 19394 17434
rect 19406 17382 19458 17434
rect 19470 17382 19522 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 2688 17323 2740 17332
rect 2688 17289 2697 17323
rect 2697 17289 2731 17323
rect 2731 17289 2740 17323
rect 2688 17280 2740 17289
rect 4620 17280 4672 17332
rect 12900 17280 12952 17332
rect 12992 17280 13044 17332
rect 11428 17212 11480 17264
rect 1400 17144 1452 17196
rect 5632 17144 5684 17196
rect 5724 17144 5776 17196
rect 6644 17144 6696 17196
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 11612 17144 11664 17196
rect 4252 17119 4304 17128
rect 4252 17085 4261 17119
rect 4261 17085 4295 17119
rect 4295 17085 4304 17119
rect 4252 17076 4304 17085
rect 4344 17119 4396 17128
rect 4344 17085 4353 17119
rect 4353 17085 4387 17119
rect 4387 17085 4396 17119
rect 4344 17076 4396 17085
rect 7656 17076 7708 17128
rect 10140 17076 10192 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 3516 16940 3568 16992
rect 5264 16940 5316 16992
rect 6184 16940 6236 16992
rect 8576 16983 8628 16992
rect 8576 16949 8585 16983
rect 8585 16949 8619 16983
rect 8619 16949 8628 16983
rect 8576 16940 8628 16949
rect 9588 16983 9640 16992
rect 9588 16949 9597 16983
rect 9597 16949 9631 16983
rect 9631 16949 9640 16983
rect 9588 16940 9640 16949
rect 12532 17144 12584 17196
rect 12624 17187 12676 17196
rect 12624 17153 12633 17187
rect 12633 17153 12667 17187
rect 12667 17153 12676 17187
rect 12624 17144 12676 17153
rect 13084 17212 13136 17264
rect 13636 17212 13688 17264
rect 17960 17212 18012 17264
rect 13912 17144 13964 17196
rect 14464 17144 14516 17196
rect 18696 17144 18748 17196
rect 19616 17144 19668 17196
rect 13544 16940 13596 16992
rect 13728 16940 13780 16992
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 18144 16940 18196 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 10214 16838 10266 16890
rect 10278 16838 10330 16890
rect 10342 16838 10394 16890
rect 10406 16838 10458 16890
rect 10470 16838 10522 16890
rect 16214 16838 16266 16890
rect 16278 16838 16330 16890
rect 16342 16838 16394 16890
rect 16406 16838 16458 16890
rect 16470 16838 16522 16890
rect 3884 16736 3936 16788
rect 6184 16779 6236 16788
rect 6184 16745 6214 16779
rect 6214 16745 6236 16779
rect 6184 16736 6236 16745
rect 7656 16779 7708 16788
rect 7656 16745 7665 16779
rect 7665 16745 7699 16779
rect 7699 16745 7708 16779
rect 7656 16736 7708 16745
rect 10140 16736 10192 16788
rect 10600 16736 10652 16788
rect 10876 16736 10928 16788
rect 13728 16736 13780 16788
rect 2044 16600 2096 16652
rect 5264 16532 5316 16584
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 14280 16600 14332 16652
rect 940 16464 992 16516
rect 2688 16464 2740 16516
rect 1676 16396 1728 16448
rect 3332 16396 3384 16448
rect 3424 16396 3476 16448
rect 3516 16396 3568 16448
rect 5080 16464 5132 16516
rect 5540 16507 5592 16516
rect 5540 16473 5558 16507
rect 5558 16473 5592 16507
rect 5540 16464 5592 16473
rect 4620 16396 4672 16448
rect 4896 16396 4948 16448
rect 6644 16464 6696 16516
rect 6828 16396 6880 16448
rect 8668 16532 8720 16584
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 11428 16575 11480 16584
rect 11428 16541 11462 16575
rect 11462 16541 11480 16575
rect 11428 16532 11480 16541
rect 14096 16532 14148 16584
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 18604 16779 18656 16788
rect 18604 16745 18613 16779
rect 18613 16745 18647 16779
rect 18647 16745 18656 16779
rect 18604 16736 18656 16745
rect 18696 16736 18748 16788
rect 19616 16736 19668 16788
rect 17316 16600 17368 16652
rect 17592 16600 17644 16652
rect 17684 16532 17736 16584
rect 17960 16532 18012 16584
rect 9680 16464 9732 16516
rect 11888 16464 11940 16516
rect 8300 16396 8352 16448
rect 8668 16396 8720 16448
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 8944 16396 8996 16405
rect 12532 16439 12584 16448
rect 12532 16405 12541 16439
rect 12541 16405 12575 16439
rect 12575 16405 12584 16439
rect 12532 16396 12584 16405
rect 17592 16507 17644 16516
rect 17592 16473 17601 16507
rect 17601 16473 17635 16507
rect 17635 16473 17644 16507
rect 17592 16464 17644 16473
rect 18052 16464 18104 16516
rect 14924 16396 14976 16448
rect 18972 16464 19024 16516
rect 19064 16507 19116 16516
rect 19064 16473 19073 16507
rect 19073 16473 19107 16507
rect 19107 16473 19116 16507
rect 19064 16464 19116 16473
rect 19708 16532 19760 16584
rect 19616 16439 19668 16448
rect 19616 16405 19625 16439
rect 19625 16405 19659 16439
rect 19659 16405 19668 16439
rect 19616 16396 19668 16405
rect 7214 16294 7266 16346
rect 7278 16294 7330 16346
rect 7342 16294 7394 16346
rect 7406 16294 7458 16346
rect 7470 16294 7522 16346
rect 13214 16294 13266 16346
rect 13278 16294 13330 16346
rect 13342 16294 13394 16346
rect 13406 16294 13458 16346
rect 13470 16294 13522 16346
rect 19214 16294 19266 16346
rect 19278 16294 19330 16346
rect 19342 16294 19394 16346
rect 19406 16294 19458 16346
rect 19470 16294 19522 16346
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 5264 16192 5316 16244
rect 5356 16192 5408 16244
rect 3424 16167 3476 16176
rect 1400 16056 1452 16108
rect 3424 16133 3433 16167
rect 3433 16133 3467 16167
rect 3467 16133 3476 16167
rect 3424 16124 3476 16133
rect 3516 16124 3568 16176
rect 8944 16192 8996 16244
rect 8852 16124 8904 16176
rect 9680 16235 9732 16244
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 15108 16192 15160 16244
rect 15476 16192 15528 16244
rect 19616 16192 19668 16244
rect 3332 16099 3384 16108
rect 3332 16065 3341 16099
rect 3341 16065 3375 16099
rect 3375 16065 3384 16099
rect 3332 16056 3384 16065
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 5080 16099 5132 16108
rect 5080 16065 5089 16099
rect 5089 16065 5123 16099
rect 5123 16065 5132 16099
rect 5080 16056 5132 16065
rect 9772 16056 9824 16108
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 3884 15988 3936 16040
rect 10140 16099 10192 16108
rect 10140 16065 10149 16099
rect 10149 16065 10183 16099
rect 10183 16065 10192 16099
rect 10140 16056 10192 16065
rect 12992 16056 13044 16108
rect 3792 15920 3844 15972
rect 12808 15988 12860 16040
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 15660 16056 15712 16108
rect 18972 16124 19024 16176
rect 19892 16124 19944 16176
rect 7932 15852 7984 15904
rect 8300 15852 8352 15904
rect 12440 15852 12492 15904
rect 14096 15852 14148 15904
rect 14372 15852 14424 15904
rect 16120 15920 16172 15972
rect 18144 16099 18196 16108
rect 18144 16065 18153 16099
rect 18153 16065 18187 16099
rect 18187 16065 18196 16099
rect 18144 16056 18196 16065
rect 15292 15852 15344 15904
rect 15384 15852 15436 15904
rect 17868 15852 17920 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 10214 15750 10266 15802
rect 10278 15750 10330 15802
rect 10342 15750 10394 15802
rect 10406 15750 10458 15802
rect 10470 15750 10522 15802
rect 16214 15750 16266 15802
rect 16278 15750 16330 15802
rect 16342 15750 16394 15802
rect 16406 15750 16458 15802
rect 16470 15750 16522 15802
rect 3516 15580 3568 15632
rect 6092 15580 6144 15632
rect 12440 15648 12492 15700
rect 12532 15648 12584 15700
rect 1676 15444 1728 15496
rect 11152 15512 11204 15564
rect 7840 15376 7892 15428
rect 8852 15376 8904 15428
rect 9864 15376 9916 15428
rect 13636 15648 13688 15700
rect 13912 15691 13964 15700
rect 13912 15657 13921 15691
rect 13921 15657 13955 15691
rect 13955 15657 13964 15691
rect 13912 15648 13964 15657
rect 14096 15648 14148 15700
rect 12992 15580 13044 15632
rect 15568 15648 15620 15700
rect 16120 15648 16172 15700
rect 18236 15580 18288 15632
rect 12716 15444 12768 15496
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 14188 15444 14240 15496
rect 14372 15487 14424 15496
rect 14372 15453 14406 15487
rect 14406 15453 14424 15487
rect 14372 15444 14424 15453
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17316 15444 17368 15453
rect 17592 15444 17644 15496
rect 17868 15444 17920 15496
rect 20260 15444 20312 15496
rect 1860 15308 1912 15360
rect 6000 15308 6052 15360
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 7012 15308 7064 15317
rect 12532 15308 12584 15360
rect 14648 15376 14700 15428
rect 17960 15376 18012 15428
rect 15660 15308 15712 15360
rect 18236 15308 18288 15360
rect 7214 15206 7266 15258
rect 7278 15206 7330 15258
rect 7342 15206 7394 15258
rect 7406 15206 7458 15258
rect 7470 15206 7522 15258
rect 13214 15206 13266 15258
rect 13278 15206 13330 15258
rect 13342 15206 13394 15258
rect 13406 15206 13458 15258
rect 13470 15206 13522 15258
rect 19214 15206 19266 15258
rect 19278 15206 19330 15258
rect 19342 15206 19394 15258
rect 19406 15206 19458 15258
rect 19470 15206 19522 15258
rect 1676 15104 1728 15156
rect 3516 15036 3568 15088
rect 3792 15079 3844 15088
rect 3792 15045 3801 15079
rect 3801 15045 3835 15079
rect 3835 15045 3844 15079
rect 3792 15036 3844 15045
rect 3884 15079 3936 15088
rect 3884 15045 3893 15079
rect 3893 15045 3927 15079
rect 3927 15045 3936 15079
rect 3884 15036 3936 15045
rect 7012 15104 7064 15156
rect 9772 15104 9824 15156
rect 3332 15011 3384 15020
rect 3332 14977 3341 15011
rect 3341 14977 3375 15011
rect 3375 14977 3384 15011
rect 3332 14968 3384 14977
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 3976 15011 4028 15020
rect 3976 14977 3985 15011
rect 3985 14977 4019 15011
rect 4019 14977 4028 15011
rect 3976 14968 4028 14977
rect 4068 14968 4120 15020
rect 7748 14968 7800 15020
rect 1768 14764 1820 14816
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 6000 14943 6052 14952
rect 6000 14909 6009 14943
rect 6009 14909 6043 14943
rect 6043 14909 6052 14943
rect 6000 14900 6052 14909
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 10600 14968 10652 14977
rect 10784 15011 10836 15020
rect 10784 14977 10793 15011
rect 10793 14977 10827 15011
rect 10827 14977 10836 15011
rect 10784 14968 10836 14977
rect 11152 14968 11204 15020
rect 11704 14968 11756 15020
rect 12716 15104 12768 15156
rect 12992 15104 13044 15156
rect 15660 15104 15712 15156
rect 19892 15147 19944 15156
rect 19892 15113 19901 15147
rect 19901 15113 19935 15147
rect 19935 15113 19944 15147
rect 19892 15104 19944 15113
rect 12532 15036 12584 15088
rect 13084 15036 13136 15088
rect 14648 15036 14700 15088
rect 19064 15036 19116 15088
rect 12440 14968 12492 15020
rect 18144 14968 18196 15020
rect 10140 14832 10192 14884
rect 14188 14943 14240 14952
rect 14188 14909 14197 14943
rect 14197 14909 14231 14943
rect 14231 14909 14240 14943
rect 14188 14900 14240 14909
rect 3148 14807 3200 14816
rect 3148 14773 3157 14807
rect 3157 14773 3191 14807
rect 3191 14773 3200 14807
rect 3148 14764 3200 14773
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 6368 14764 6420 14816
rect 7656 14764 7708 14816
rect 8944 14807 8996 14816
rect 8944 14773 8953 14807
rect 8953 14773 8987 14807
rect 8987 14773 8996 14807
rect 8944 14764 8996 14773
rect 9680 14807 9732 14816
rect 9680 14773 9689 14807
rect 9689 14773 9723 14807
rect 9723 14773 9732 14807
rect 9680 14764 9732 14773
rect 10048 14764 10100 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 10214 14662 10266 14714
rect 10278 14662 10330 14714
rect 10342 14662 10394 14714
rect 10406 14662 10458 14714
rect 10470 14662 10522 14714
rect 16214 14662 16266 14714
rect 16278 14662 16330 14714
rect 16342 14662 16394 14714
rect 16406 14662 16458 14714
rect 16470 14662 16522 14714
rect 1676 14560 1728 14612
rect 3148 14560 3200 14612
rect 3976 14560 4028 14612
rect 10784 14603 10836 14612
rect 10784 14569 10793 14603
rect 10793 14569 10827 14603
rect 10827 14569 10836 14603
rect 10784 14560 10836 14569
rect 12440 14560 12492 14612
rect 17408 14560 17460 14612
rect 7656 14424 7708 14476
rect 7932 14424 7984 14476
rect 8944 14424 8996 14476
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 14188 14424 14240 14476
rect 15292 14467 15344 14476
rect 15292 14433 15301 14467
rect 15301 14433 15335 14467
rect 15335 14433 15344 14467
rect 15292 14424 15344 14433
rect 16672 14424 16724 14476
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 1860 14399 1912 14408
rect 1860 14365 1869 14399
rect 1869 14365 1903 14399
rect 1903 14365 1912 14399
rect 1860 14356 1912 14365
rect 5816 14356 5868 14408
rect 10600 14356 10652 14408
rect 12532 14399 12584 14408
rect 12532 14365 12550 14399
rect 12550 14365 12584 14399
rect 12532 14356 12584 14365
rect 17132 14399 17184 14408
rect 17132 14365 17134 14399
rect 17134 14365 17168 14399
rect 17168 14365 17184 14399
rect 17132 14356 17184 14365
rect 4068 14288 4120 14340
rect 5172 14331 5224 14340
rect 5172 14297 5181 14331
rect 5181 14297 5215 14331
rect 5215 14297 5224 14331
rect 5172 14288 5224 14297
rect 6920 14331 6972 14340
rect 6920 14297 6929 14331
rect 6929 14297 6963 14331
rect 6963 14297 6972 14331
rect 6920 14288 6972 14297
rect 7748 14288 7800 14340
rect 9312 14331 9364 14340
rect 9312 14297 9321 14331
rect 9321 14297 9355 14331
rect 9355 14297 9364 14331
rect 9312 14288 9364 14297
rect 9864 14288 9916 14340
rect 15660 14288 15712 14340
rect 18144 14356 18196 14408
rect 7656 14220 7708 14272
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 17316 14263 17368 14272
rect 17316 14229 17325 14263
rect 17325 14229 17359 14263
rect 17359 14229 17368 14263
rect 17316 14220 17368 14229
rect 18972 14263 19024 14272
rect 18972 14229 18981 14263
rect 18981 14229 19015 14263
rect 19015 14229 19024 14263
rect 18972 14220 19024 14229
rect 7214 14118 7266 14170
rect 7278 14118 7330 14170
rect 7342 14118 7394 14170
rect 7406 14118 7458 14170
rect 7470 14118 7522 14170
rect 13214 14118 13266 14170
rect 13278 14118 13330 14170
rect 13342 14118 13394 14170
rect 13406 14118 13458 14170
rect 13470 14118 13522 14170
rect 19214 14118 19266 14170
rect 19278 14118 19330 14170
rect 19342 14118 19394 14170
rect 19406 14118 19458 14170
rect 19470 14118 19522 14170
rect 3332 14016 3384 14068
rect 3976 14016 4028 14068
rect 5724 14016 5776 14068
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 3516 13948 3568 14000
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 4068 13812 4120 13864
rect 5632 13880 5684 13932
rect 6368 14016 6420 14068
rect 6092 13880 6144 13932
rect 5356 13812 5408 13864
rect 6920 13948 6972 14000
rect 7656 14059 7708 14068
rect 7656 14025 7665 14059
rect 7665 14025 7699 14059
rect 7699 14025 7708 14059
rect 7656 14016 7708 14025
rect 7840 13948 7892 14000
rect 9312 14016 9364 14068
rect 11704 14016 11756 14068
rect 12808 14016 12860 14068
rect 16580 14016 16632 14068
rect 18144 14059 18196 14068
rect 18144 14025 18153 14059
rect 18153 14025 18187 14059
rect 18187 14025 18196 14059
rect 18144 14016 18196 14025
rect 9680 13948 9732 14000
rect 14556 13991 14608 14000
rect 14556 13957 14565 13991
rect 14565 13957 14599 13991
rect 14599 13957 14608 13991
rect 14556 13948 14608 13957
rect 8760 13880 8812 13932
rect 15752 13880 15804 13932
rect 18972 13948 19024 14000
rect 18052 13812 18104 13864
rect 1584 13744 1636 13796
rect 2688 13744 2740 13796
rect 10048 13744 10100 13796
rect 6000 13719 6052 13728
rect 6000 13685 6009 13719
rect 6009 13685 6043 13719
rect 6043 13685 6052 13719
rect 6000 13676 6052 13685
rect 8300 13719 8352 13728
rect 8300 13685 8309 13719
rect 8309 13685 8343 13719
rect 8343 13685 8352 13719
rect 8300 13676 8352 13685
rect 10600 13676 10652 13728
rect 16580 13676 16632 13728
rect 17132 13676 17184 13728
rect 19984 13719 20036 13728
rect 19984 13685 19993 13719
rect 19993 13685 20027 13719
rect 20027 13685 20036 13719
rect 19984 13676 20036 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 10214 13574 10266 13626
rect 10278 13574 10330 13626
rect 10342 13574 10394 13626
rect 10406 13574 10458 13626
rect 10470 13574 10522 13626
rect 16214 13574 16266 13626
rect 16278 13574 16330 13626
rect 16342 13574 16394 13626
rect 16406 13574 16458 13626
rect 16470 13574 16522 13626
rect 6000 13472 6052 13524
rect 7840 13472 7892 13524
rect 4528 13379 4580 13388
rect 4528 13345 4537 13379
rect 4537 13345 4571 13379
rect 4571 13345 4580 13379
rect 4528 13336 4580 13345
rect 5448 13336 5500 13388
rect 9680 13336 9732 13388
rect 9956 13336 10008 13388
rect 2688 13268 2740 13320
rect 3516 13311 3568 13320
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 7748 13268 7800 13320
rect 9496 13268 9548 13320
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 2504 13175 2556 13184
rect 2504 13141 2513 13175
rect 2513 13141 2547 13175
rect 2547 13141 2556 13175
rect 2504 13132 2556 13141
rect 3148 13132 3200 13184
rect 4160 13175 4212 13184
rect 4160 13141 4169 13175
rect 4169 13141 4203 13175
rect 4203 13141 4212 13175
rect 4160 13132 4212 13141
rect 4344 13175 4396 13184
rect 4344 13141 4353 13175
rect 4353 13141 4387 13175
rect 4387 13141 4396 13175
rect 4344 13132 4396 13141
rect 6920 13132 6972 13184
rect 9312 13243 9364 13252
rect 9312 13209 9321 13243
rect 9321 13209 9355 13243
rect 9355 13209 9364 13243
rect 9312 13200 9364 13209
rect 9772 13200 9824 13252
rect 10600 13336 10652 13388
rect 17040 13472 17092 13524
rect 17408 13472 17460 13524
rect 17868 13472 17920 13524
rect 15660 13447 15712 13456
rect 15660 13413 15669 13447
rect 15669 13413 15703 13447
rect 15703 13413 15712 13447
rect 15660 13404 15712 13413
rect 16580 13404 16632 13456
rect 14188 13336 14240 13388
rect 8944 13175 8996 13184
rect 8944 13141 8953 13175
rect 8953 13141 8987 13175
rect 8987 13141 8996 13175
rect 8944 13132 8996 13141
rect 10876 13200 10928 13252
rect 12164 13243 12216 13252
rect 12164 13209 12173 13243
rect 12173 13209 12207 13243
rect 12207 13209 12216 13243
rect 12164 13200 12216 13209
rect 14556 13243 14608 13252
rect 14556 13209 14579 13243
rect 14579 13209 14608 13243
rect 14556 13200 14608 13209
rect 12072 13175 12124 13184
rect 12072 13141 12081 13175
rect 12081 13141 12115 13175
rect 12115 13141 12124 13175
rect 12072 13132 12124 13141
rect 13084 13132 13136 13184
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 13728 13175 13780 13184
rect 13728 13141 13737 13175
rect 13737 13141 13771 13175
rect 13771 13141 13780 13175
rect 13728 13132 13780 13141
rect 16580 13268 16632 13320
rect 17684 13268 17736 13320
rect 18052 13268 18104 13320
rect 16028 13132 16080 13184
rect 16304 13175 16356 13184
rect 16304 13141 16313 13175
rect 16313 13141 16347 13175
rect 16347 13141 16356 13175
rect 16304 13132 16356 13141
rect 16672 13132 16724 13184
rect 7214 13030 7266 13082
rect 7278 13030 7330 13082
rect 7342 13030 7394 13082
rect 7406 13030 7458 13082
rect 7470 13030 7522 13082
rect 13214 13030 13266 13082
rect 13278 13030 13330 13082
rect 13342 13030 13394 13082
rect 13406 13030 13458 13082
rect 13470 13030 13522 13082
rect 19214 13030 19266 13082
rect 19278 13030 19330 13082
rect 19342 13030 19394 13082
rect 19406 13030 19458 13082
rect 19470 13030 19522 13082
rect 2688 12928 2740 12980
rect 3148 12928 3200 12980
rect 4344 12928 4396 12980
rect 6368 12928 6420 12980
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 9128 12928 9180 12980
rect 1400 12724 1452 12776
rect 1676 12656 1728 12708
rect 2504 12792 2556 12844
rect 3976 12792 4028 12844
rect 5724 12792 5776 12844
rect 7104 12860 7156 12912
rect 1768 12631 1820 12640
rect 1768 12597 1777 12631
rect 1777 12597 1811 12631
rect 1811 12597 1820 12631
rect 1768 12588 1820 12597
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 1952 12588 2004 12597
rect 3424 12724 3476 12776
rect 5448 12724 5500 12776
rect 9404 12792 9456 12844
rect 9864 12928 9916 12980
rect 10876 12928 10928 12980
rect 12072 12928 12124 12980
rect 13636 12928 13688 12980
rect 14096 12928 14148 12980
rect 14556 12928 14608 12980
rect 9956 12860 10008 12912
rect 15292 12903 15344 12912
rect 15292 12869 15310 12903
rect 15310 12869 15344 12903
rect 15292 12860 15344 12869
rect 8392 12724 8444 12776
rect 9496 12724 9548 12776
rect 9772 12724 9824 12776
rect 4712 12588 4764 12640
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 13084 12792 13136 12844
rect 16028 12928 16080 12980
rect 16672 12928 16724 12980
rect 17132 12928 17184 12980
rect 19248 12928 19300 12980
rect 16304 12860 16356 12912
rect 17868 12903 17920 12912
rect 17868 12869 17886 12903
rect 17886 12869 17920 12903
rect 17868 12860 17920 12869
rect 18512 12903 18564 12912
rect 18512 12869 18521 12903
rect 18521 12869 18555 12903
rect 18555 12869 18564 12903
rect 18512 12860 18564 12869
rect 18972 12860 19024 12912
rect 19984 12860 20036 12912
rect 18052 12792 18104 12844
rect 13636 12767 13688 12776
rect 13636 12733 13645 12767
rect 13645 12733 13679 12767
rect 13679 12733 13688 12767
rect 13636 12724 13688 12733
rect 15568 12767 15620 12776
rect 15568 12733 15577 12767
rect 15577 12733 15611 12767
rect 15611 12733 15620 12767
rect 15568 12724 15620 12733
rect 19524 12792 19576 12844
rect 18788 12724 18840 12776
rect 15660 12656 15712 12708
rect 10140 12588 10192 12597
rect 13728 12588 13780 12640
rect 15292 12588 15344 12640
rect 17132 12656 17184 12708
rect 18880 12699 18932 12708
rect 18880 12665 18889 12699
rect 18889 12665 18923 12699
rect 18923 12665 18932 12699
rect 18880 12656 18932 12665
rect 18328 12631 18380 12640
rect 18328 12597 18337 12631
rect 18337 12597 18371 12631
rect 18371 12597 18380 12631
rect 18328 12588 18380 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 10214 12486 10266 12538
rect 10278 12486 10330 12538
rect 10342 12486 10394 12538
rect 10406 12486 10458 12538
rect 10470 12486 10522 12538
rect 16214 12486 16266 12538
rect 16278 12486 16330 12538
rect 16342 12486 16394 12538
rect 16406 12486 16458 12538
rect 16470 12486 16522 12538
rect 1952 12384 2004 12436
rect 3516 12384 3568 12436
rect 5356 12384 5408 12436
rect 8392 12384 8444 12436
rect 9312 12427 9364 12436
rect 9312 12393 9321 12427
rect 9321 12393 9355 12427
rect 9355 12393 9364 12427
rect 9312 12384 9364 12393
rect 13728 12384 13780 12436
rect 19248 12427 19300 12436
rect 19248 12393 19257 12427
rect 19257 12393 19291 12427
rect 19291 12393 19300 12427
rect 19248 12384 19300 12393
rect 18604 12316 18656 12368
rect 19524 12316 19576 12368
rect 1400 12180 1452 12232
rect 2596 12248 2648 12300
rect 1860 12223 1912 12232
rect 1860 12189 1869 12223
rect 1869 12189 1903 12223
rect 1903 12189 1912 12223
rect 1860 12180 1912 12189
rect 3240 12180 3292 12232
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 2412 12112 2464 12164
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 4712 12180 4764 12232
rect 8760 12223 8812 12232
rect 8760 12189 8769 12223
rect 8769 12189 8803 12223
rect 8803 12189 8812 12223
rect 8760 12180 8812 12189
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9588 12223 9640 12232
rect 9588 12189 9597 12223
rect 9597 12189 9631 12223
rect 9631 12189 9640 12223
rect 9588 12180 9640 12189
rect 10140 12180 10192 12232
rect 12716 12180 12768 12232
rect 14096 12180 14148 12232
rect 14372 12180 14424 12232
rect 15568 12223 15620 12232
rect 15568 12189 15577 12223
rect 15577 12189 15611 12223
rect 15611 12189 15620 12223
rect 15568 12180 15620 12189
rect 18880 12248 18932 12300
rect 18696 12180 18748 12232
rect 3516 12112 3568 12164
rect 4068 12155 4120 12164
rect 4068 12121 4077 12155
rect 4077 12121 4111 12155
rect 4111 12121 4120 12155
rect 4068 12112 4120 12121
rect 5264 12112 5316 12164
rect 15936 12155 15988 12164
rect 15936 12121 15970 12155
rect 15970 12121 15988 12155
rect 12532 12044 12584 12096
rect 15936 12112 15988 12121
rect 18052 12112 18104 12164
rect 20168 12155 20220 12164
rect 20168 12121 20177 12155
rect 20177 12121 20211 12155
rect 20211 12121 20220 12155
rect 20168 12112 20220 12121
rect 15660 12044 15712 12096
rect 16672 12044 16724 12096
rect 18144 12044 18196 12096
rect 19892 12087 19944 12096
rect 19892 12053 19901 12087
rect 19901 12053 19935 12087
rect 19935 12053 19944 12087
rect 19892 12044 19944 12053
rect 7214 11942 7266 11994
rect 7278 11942 7330 11994
rect 7342 11942 7394 11994
rect 7406 11942 7458 11994
rect 7470 11942 7522 11994
rect 13214 11942 13266 11994
rect 13278 11942 13330 11994
rect 13342 11942 13394 11994
rect 13406 11942 13458 11994
rect 13470 11942 13522 11994
rect 19214 11942 19266 11994
rect 19278 11942 19330 11994
rect 19342 11942 19394 11994
rect 19406 11942 19458 11994
rect 19470 11942 19522 11994
rect 1584 11840 1636 11892
rect 2412 11840 2464 11892
rect 4068 11840 4120 11892
rect 13084 11840 13136 11892
rect 13636 11840 13688 11892
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 3424 11704 3476 11756
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 14372 11772 14424 11824
rect 6828 11636 6880 11688
rect 8944 11636 8996 11688
rect 11152 11636 11204 11688
rect 15752 11704 15804 11756
rect 15936 11772 15988 11824
rect 16764 11840 16816 11892
rect 18052 11840 18104 11892
rect 17960 11815 18012 11824
rect 17960 11781 17969 11815
rect 17969 11781 18003 11815
rect 18003 11781 18012 11815
rect 17960 11772 18012 11781
rect 17316 11704 17368 11756
rect 19892 11840 19944 11892
rect 18604 11772 18656 11824
rect 19064 11772 19116 11824
rect 20168 11772 20220 11824
rect 18328 11704 18380 11756
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 16764 11568 16816 11620
rect 8392 11500 8444 11552
rect 9864 11500 9916 11552
rect 10876 11500 10928 11552
rect 14372 11500 14424 11552
rect 16672 11500 16724 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 17132 11543 17184 11552
rect 17132 11509 17141 11543
rect 17141 11509 17175 11543
rect 17175 11509 17184 11543
rect 17132 11500 17184 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 10214 11398 10266 11450
rect 10278 11398 10330 11450
rect 10342 11398 10394 11450
rect 10406 11398 10458 11450
rect 10470 11398 10522 11450
rect 16214 11398 16266 11450
rect 16278 11398 16330 11450
rect 16342 11398 16394 11450
rect 16406 11398 16458 11450
rect 16470 11398 16522 11450
rect 1676 11296 1728 11348
rect 5264 11296 5316 11348
rect 7932 11296 7984 11348
rect 9772 11296 9824 11348
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 17224 11296 17276 11348
rect 17592 11339 17644 11348
rect 17592 11305 17601 11339
rect 17601 11305 17635 11339
rect 17635 11305 17644 11339
rect 17592 11296 17644 11305
rect 18052 11296 18104 11348
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 9036 11228 9088 11280
rect 5264 11203 5316 11212
rect 5264 11169 5273 11203
rect 5273 11169 5307 11203
rect 5307 11169 5316 11203
rect 5264 11160 5316 11169
rect 8944 11160 8996 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 6920 11092 6972 11144
rect 10600 11160 10652 11212
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 7012 10999 7064 11008
rect 7012 10965 7021 10999
rect 7021 10965 7055 10999
rect 7055 10965 7064 10999
rect 7012 10956 7064 10965
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 8208 11067 8260 11076
rect 8208 11033 8217 11067
rect 8217 11033 8251 11067
rect 8251 11033 8260 11067
rect 8208 11024 8260 11033
rect 8484 11024 8536 11076
rect 9404 11024 9456 11076
rect 11060 11024 11112 11076
rect 8116 10999 8168 11008
rect 8116 10965 8125 10999
rect 8125 10965 8159 10999
rect 8159 10965 8168 10999
rect 8116 10956 8168 10965
rect 13912 11160 13964 11212
rect 17776 11160 17828 11212
rect 15936 11092 15988 11144
rect 13820 11024 13872 11076
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 13084 10956 13136 11008
rect 15844 11024 15896 11076
rect 16764 11024 16816 11076
rect 19800 11092 19852 11144
rect 19708 11067 19760 11076
rect 19708 11033 19717 11067
rect 19717 11033 19751 11067
rect 19751 11033 19760 11067
rect 19708 11024 19760 11033
rect 20076 10956 20128 11008
rect 7214 10854 7266 10906
rect 7278 10854 7330 10906
rect 7342 10854 7394 10906
rect 7406 10854 7458 10906
rect 7470 10854 7522 10906
rect 13214 10854 13266 10906
rect 13278 10854 13330 10906
rect 13342 10854 13394 10906
rect 13406 10854 13458 10906
rect 13470 10854 13522 10906
rect 19214 10854 19266 10906
rect 19278 10854 19330 10906
rect 19342 10854 19394 10906
rect 19406 10854 19458 10906
rect 19470 10854 19522 10906
rect 4620 10752 4672 10804
rect 4804 10752 4856 10804
rect 5172 10684 5224 10736
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 7104 10752 7156 10804
rect 7656 10752 7708 10804
rect 9036 10752 9088 10804
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 4804 10659 4856 10668
rect 4804 10625 4813 10659
rect 4813 10625 4847 10659
rect 4847 10625 4856 10659
rect 4804 10616 4856 10625
rect 5540 10616 5592 10668
rect 4896 10591 4948 10600
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 7012 10659 7064 10668
rect 7012 10625 7021 10659
rect 7021 10625 7055 10659
rect 7055 10625 7064 10659
rect 7012 10616 7064 10625
rect 6736 10548 6788 10600
rect 7472 10616 7524 10668
rect 9404 10684 9456 10736
rect 7564 10480 7616 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 7104 10455 7156 10464
rect 7104 10421 7113 10455
rect 7113 10421 7147 10455
rect 7147 10421 7156 10455
rect 7104 10412 7156 10421
rect 8024 10616 8076 10668
rect 16764 10795 16816 10804
rect 16764 10761 16773 10795
rect 16773 10761 16807 10795
rect 16807 10761 16816 10795
rect 16764 10752 16816 10761
rect 11336 10684 11388 10736
rect 12624 10684 12676 10736
rect 15200 10684 15252 10736
rect 19616 10752 19668 10804
rect 10140 10616 10192 10668
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 10876 10659 10928 10668
rect 10876 10625 10885 10659
rect 10885 10625 10919 10659
rect 10919 10625 10928 10659
rect 10876 10616 10928 10625
rect 11152 10659 11204 10668
rect 11152 10625 11155 10659
rect 11155 10625 11204 10659
rect 11152 10616 11204 10625
rect 7748 10591 7800 10600
rect 7748 10557 7757 10591
rect 7757 10557 7791 10591
rect 7791 10557 7800 10591
rect 7748 10548 7800 10557
rect 7932 10548 7984 10600
rect 8392 10548 8444 10600
rect 12440 10616 12492 10668
rect 13820 10616 13872 10668
rect 17868 10659 17920 10668
rect 17868 10625 17886 10659
rect 17886 10625 17920 10659
rect 17868 10616 17920 10625
rect 18052 10616 18104 10668
rect 18788 10616 18840 10668
rect 19708 10616 19760 10668
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 12164 10548 12216 10600
rect 14188 10591 14240 10600
rect 14188 10557 14197 10591
rect 14197 10557 14231 10591
rect 14231 10557 14240 10591
rect 14188 10548 14240 10557
rect 9864 10480 9916 10532
rect 19800 10523 19852 10532
rect 19800 10489 19809 10523
rect 19809 10489 19843 10523
rect 19843 10489 19852 10523
rect 19800 10480 19852 10489
rect 9680 10455 9732 10464
rect 9680 10421 9689 10455
rect 9689 10421 9723 10455
rect 9723 10421 9732 10455
rect 9680 10412 9732 10421
rect 9956 10412 10008 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 10784 10412 10836 10464
rect 11060 10412 11112 10464
rect 13084 10412 13136 10464
rect 19616 10455 19668 10464
rect 19616 10421 19625 10455
rect 19625 10421 19659 10455
rect 19659 10421 19668 10455
rect 19616 10412 19668 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 10214 10310 10266 10362
rect 10278 10310 10330 10362
rect 10342 10310 10394 10362
rect 10406 10310 10458 10362
rect 10470 10310 10522 10362
rect 16214 10310 16266 10362
rect 16278 10310 16330 10362
rect 16342 10310 16394 10362
rect 16406 10310 16458 10362
rect 16470 10310 16522 10362
rect 4804 10208 4856 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 7012 10208 7064 10260
rect 7748 10208 7800 10260
rect 8024 10208 8076 10260
rect 8668 10208 8720 10260
rect 9680 10208 9732 10260
rect 9772 10208 9824 10260
rect 10048 10208 10100 10260
rect 10600 10208 10652 10260
rect 14188 10208 14240 10260
rect 15936 10208 15988 10260
rect 18236 10208 18288 10260
rect 20168 10208 20220 10260
rect 7472 10072 7524 10124
rect 7748 10072 7800 10124
rect 3424 9936 3476 9988
rect 8116 10004 8168 10056
rect 10876 10072 10928 10124
rect 2780 9868 2832 9920
rect 3976 9936 4028 9988
rect 4344 9936 4396 9988
rect 6920 9936 6972 9988
rect 8760 9936 8812 9988
rect 9128 9979 9180 9988
rect 9128 9945 9137 9979
rect 9137 9945 9171 9979
rect 9171 9945 9180 9979
rect 9128 9936 9180 9945
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 6644 9868 6696 9920
rect 8024 9868 8076 9920
rect 10600 10004 10652 10056
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 9956 9936 10008 9988
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 13820 10047 13872 10056
rect 13820 10013 13829 10047
rect 13829 10013 13863 10047
rect 13863 10013 13872 10047
rect 13820 10004 13872 10013
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 16120 10004 16172 10056
rect 19616 10140 19668 10192
rect 18328 10004 18380 10056
rect 18696 10047 18748 10056
rect 18696 10013 18705 10047
rect 18705 10013 18739 10047
rect 18739 10013 18748 10047
rect 18696 10004 18748 10013
rect 14648 9979 14700 9988
rect 14648 9945 14682 9979
rect 14682 9945 14700 9979
rect 14648 9936 14700 9945
rect 10048 9868 10100 9920
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 18144 9868 18196 9877
rect 18236 9868 18288 9920
rect 20168 10004 20220 10056
rect 20812 10004 20864 10056
rect 7214 9766 7266 9818
rect 7278 9766 7330 9818
rect 7342 9766 7394 9818
rect 7406 9766 7458 9818
rect 7470 9766 7522 9818
rect 13214 9766 13266 9818
rect 13278 9766 13330 9818
rect 13342 9766 13394 9818
rect 13406 9766 13458 9818
rect 13470 9766 13522 9818
rect 19214 9766 19266 9818
rect 19278 9766 19330 9818
rect 19342 9766 19394 9818
rect 19406 9766 19458 9818
rect 19470 9766 19522 9818
rect 2780 9707 2832 9716
rect 2780 9673 2789 9707
rect 2789 9673 2823 9707
rect 2823 9673 2832 9707
rect 2780 9664 2832 9673
rect 4344 9664 4396 9716
rect 4896 9664 4948 9716
rect 5080 9664 5132 9716
rect 5632 9664 5684 9716
rect 1584 9528 1636 9580
rect 6828 9664 6880 9716
rect 6920 9707 6972 9716
rect 6920 9673 6929 9707
rect 6929 9673 6963 9707
rect 6963 9673 6972 9707
rect 6920 9664 6972 9673
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 5080 9571 5132 9580
rect 7104 9596 7156 9648
rect 5080 9537 5115 9571
rect 5115 9537 5132 9571
rect 5080 9528 5132 9537
rect 5908 9571 5960 9580
rect 5908 9537 5917 9571
rect 5917 9537 5951 9571
rect 5951 9537 5960 9571
rect 5908 9528 5960 9537
rect 1768 9367 1820 9376
rect 1768 9333 1777 9367
rect 1777 9333 1811 9367
rect 1811 9333 1820 9367
rect 1768 9324 1820 9333
rect 3976 9324 4028 9376
rect 5724 9503 5776 9512
rect 5724 9469 5733 9503
rect 5733 9469 5767 9503
rect 5767 9469 5776 9503
rect 5724 9460 5776 9469
rect 5816 9460 5868 9512
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 7104 9460 7156 9512
rect 4804 9392 4856 9444
rect 5356 9392 5408 9444
rect 4620 9324 4672 9376
rect 5080 9324 5132 9376
rect 5448 9324 5500 9376
rect 5632 9324 5684 9376
rect 6644 9392 6696 9444
rect 6736 9392 6788 9444
rect 7564 9664 7616 9716
rect 9772 9664 9824 9716
rect 9864 9664 9916 9716
rect 10784 9664 10836 9716
rect 12440 9707 12492 9716
rect 12440 9673 12449 9707
rect 12449 9673 12483 9707
rect 12483 9673 12492 9707
rect 12440 9664 12492 9673
rect 14648 9596 14700 9648
rect 18236 9664 18288 9716
rect 18788 9707 18840 9716
rect 18788 9673 18797 9707
rect 18797 9673 18831 9707
rect 18831 9673 18840 9707
rect 18788 9664 18840 9673
rect 7932 9528 7984 9580
rect 9036 9528 9088 9580
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 8208 9460 8260 9512
rect 9588 9571 9640 9580
rect 9588 9537 9597 9571
rect 9597 9537 9631 9571
rect 9631 9537 9640 9571
rect 9588 9528 9640 9537
rect 10140 9528 10192 9580
rect 12532 9528 12584 9580
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 14372 9528 14424 9580
rect 7932 9392 7984 9444
rect 9036 9392 9088 9444
rect 9312 9392 9364 9444
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8576 9324 8628 9376
rect 9220 9324 9272 9376
rect 11244 9324 11296 9376
rect 11612 9324 11664 9376
rect 15200 9324 15252 9376
rect 16580 9324 16632 9376
rect 19708 9528 19760 9580
rect 18972 9503 19024 9512
rect 18972 9469 18981 9503
rect 18981 9469 19015 9503
rect 19015 9469 19024 9503
rect 18972 9460 19024 9469
rect 20076 9324 20128 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 10214 9222 10266 9274
rect 10278 9222 10330 9274
rect 10342 9222 10394 9274
rect 10406 9222 10458 9274
rect 10470 9222 10522 9274
rect 16214 9222 16266 9274
rect 16278 9222 16330 9274
rect 16342 9222 16394 9274
rect 16406 9222 16458 9274
rect 16470 9222 16522 9274
rect 1768 9120 1820 9172
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 5632 8984 5684 9036
rect 5172 8916 5224 8968
rect 5816 9120 5868 9172
rect 5908 9120 5960 9172
rect 7012 9120 7064 9172
rect 7104 9120 7156 9172
rect 7748 9120 7800 9172
rect 9128 9120 9180 9172
rect 9220 9163 9272 9172
rect 9220 9129 9229 9163
rect 9229 9129 9263 9163
rect 9263 9129 9272 9163
rect 9220 9120 9272 9129
rect 17776 9163 17828 9172
rect 17776 9129 17785 9163
rect 17785 9129 17819 9163
rect 17819 9129 17828 9163
rect 17776 9120 17828 9129
rect 18144 9120 18196 9172
rect 4620 8848 4672 8900
rect 5356 8891 5408 8900
rect 5356 8857 5365 8891
rect 5365 8857 5399 8891
rect 5399 8857 5408 8891
rect 5356 8848 5408 8857
rect 6276 8916 6328 8968
rect 7932 8916 7984 8968
rect 8208 8916 8260 8968
rect 18052 9052 18104 9104
rect 10140 8984 10192 9036
rect 10508 8984 10560 9036
rect 11060 8984 11112 9036
rect 12440 8984 12492 9036
rect 9404 8916 9456 8968
rect 11796 8916 11848 8968
rect 16580 8984 16632 9036
rect 18144 8984 18196 9036
rect 17684 8916 17736 8968
rect 18696 9120 18748 9172
rect 7564 8848 7616 8900
rect 8760 8848 8812 8900
rect 2228 8823 2280 8832
rect 2228 8789 2237 8823
rect 2237 8789 2271 8823
rect 2271 8789 2280 8823
rect 2228 8780 2280 8789
rect 4252 8780 4304 8832
rect 4712 8780 4764 8832
rect 5264 8780 5316 8832
rect 5448 8780 5500 8832
rect 6460 8780 6512 8832
rect 7840 8780 7892 8832
rect 8024 8780 8076 8832
rect 9036 8823 9088 8832
rect 9036 8789 9045 8823
rect 9045 8789 9079 8823
rect 9079 8789 9088 8823
rect 9036 8780 9088 8789
rect 9772 8891 9824 8900
rect 9772 8857 9781 8891
rect 9781 8857 9815 8891
rect 9815 8857 9824 8891
rect 9772 8848 9824 8857
rect 10784 8848 10836 8900
rect 11336 8891 11388 8900
rect 11336 8857 11345 8891
rect 11345 8857 11379 8891
rect 11379 8857 11388 8891
rect 11336 8848 11388 8857
rect 12164 8848 12216 8900
rect 17592 8891 17644 8900
rect 17592 8857 17601 8891
rect 17601 8857 17635 8891
rect 17635 8857 17644 8891
rect 17592 8848 17644 8857
rect 11152 8780 11204 8832
rect 12072 8780 12124 8832
rect 12808 8780 12860 8832
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 15384 8780 15436 8832
rect 17316 8780 17368 8832
rect 18052 8891 18104 8900
rect 18052 8857 18061 8891
rect 18061 8857 18095 8891
rect 18095 8857 18104 8891
rect 18052 8848 18104 8857
rect 18788 8780 18840 8832
rect 7214 8678 7266 8730
rect 7278 8678 7330 8730
rect 7342 8678 7394 8730
rect 7406 8678 7458 8730
rect 7470 8678 7522 8730
rect 13214 8678 13266 8730
rect 13278 8678 13330 8730
rect 13342 8678 13394 8730
rect 13406 8678 13458 8730
rect 13470 8678 13522 8730
rect 19214 8678 19266 8730
rect 19278 8678 19330 8730
rect 19342 8678 19394 8730
rect 19406 8678 19458 8730
rect 19470 8678 19522 8730
rect 2228 8576 2280 8628
rect 5264 8576 5316 8628
rect 5816 8576 5868 8628
rect 7012 8576 7064 8628
rect 4252 8551 4304 8560
rect 4252 8517 4261 8551
rect 4261 8517 4295 8551
rect 4295 8517 4304 8551
rect 4252 8508 4304 8517
rect 4436 8551 4488 8560
rect 4436 8517 4471 8551
rect 4471 8517 4488 8551
rect 4436 8508 4488 8517
rect 4712 8551 4764 8560
rect 4712 8517 4721 8551
rect 4721 8517 4755 8551
rect 4755 8517 4764 8551
rect 4712 8508 4764 8517
rect 6920 8551 6972 8560
rect 6920 8517 6929 8551
rect 6929 8517 6963 8551
rect 6963 8517 6972 8551
rect 6920 8508 6972 8517
rect 4620 8415 4672 8424
rect 4620 8381 4629 8415
rect 4629 8381 4663 8415
rect 4663 8381 4672 8415
rect 4620 8372 4672 8381
rect 5172 8483 5224 8492
rect 5172 8449 5178 8483
rect 5178 8449 5212 8483
rect 5212 8449 5224 8483
rect 5172 8440 5224 8449
rect 5632 8440 5684 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 5908 8440 5960 8492
rect 6644 8440 6696 8492
rect 8208 8508 8260 8560
rect 8760 8508 8812 8560
rect 9312 8576 9364 8628
rect 9404 8508 9456 8560
rect 10508 8508 10560 8560
rect 12624 8576 12676 8628
rect 12808 8576 12860 8628
rect 13544 8576 13596 8628
rect 5632 8304 5684 8356
rect 6276 8304 6328 8356
rect 6736 8304 6788 8356
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 10968 8483 11020 8492
rect 10968 8449 10977 8483
rect 10977 8449 11011 8483
rect 11011 8449 11020 8483
rect 10968 8440 11020 8449
rect 12440 8508 12492 8560
rect 13544 8440 13596 8492
rect 14280 8576 14332 8628
rect 18052 8576 18104 8628
rect 18972 8576 19024 8628
rect 19708 8576 19760 8628
rect 15936 8508 15988 8560
rect 16580 8508 16632 8560
rect 15844 8440 15896 8492
rect 17684 8440 17736 8492
rect 19064 8440 19116 8492
rect 11428 8372 11480 8424
rect 11612 8415 11664 8424
rect 11612 8381 11621 8415
rect 11621 8381 11655 8415
rect 11655 8381 11664 8415
rect 11612 8372 11664 8381
rect 1768 8279 1820 8288
rect 1768 8245 1777 8279
rect 1777 8245 1811 8279
rect 1811 8245 1820 8279
rect 1768 8236 1820 8245
rect 2964 8236 3016 8288
rect 4896 8236 4948 8288
rect 5172 8236 5224 8288
rect 6368 8279 6420 8288
rect 6368 8245 6377 8279
rect 6377 8245 6411 8279
rect 6411 8245 6420 8279
rect 6368 8236 6420 8245
rect 6644 8236 6696 8288
rect 7472 8279 7524 8288
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 8392 8236 8444 8288
rect 10140 8304 10192 8356
rect 13820 8372 13872 8424
rect 15568 8304 15620 8356
rect 9864 8236 9916 8288
rect 12256 8236 12308 8288
rect 13084 8236 13136 8288
rect 15384 8236 15436 8288
rect 16028 8236 16080 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 10214 8134 10266 8186
rect 10278 8134 10330 8186
rect 10342 8134 10394 8186
rect 10406 8134 10458 8186
rect 10470 8134 10522 8186
rect 16214 8134 16266 8186
rect 16278 8134 16330 8186
rect 16342 8134 16394 8186
rect 16406 8134 16458 8186
rect 16470 8134 16522 8186
rect 3608 8032 3660 8084
rect 5816 8032 5868 8084
rect 5632 7964 5684 8016
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 2504 7803 2556 7812
rect 2504 7769 2513 7803
rect 2513 7769 2547 7803
rect 2547 7769 2556 7803
rect 2504 7760 2556 7769
rect 5448 7828 5500 7880
rect 6460 8007 6512 8016
rect 6460 7973 6469 8007
rect 6469 7973 6503 8007
rect 6503 7973 6512 8007
rect 6460 7964 6512 7973
rect 10600 8032 10652 8084
rect 10784 8075 10836 8084
rect 10784 8041 10793 8075
rect 10793 8041 10827 8075
rect 10827 8041 10836 8075
rect 10784 8032 10836 8041
rect 16028 8032 16080 8084
rect 17224 8075 17276 8084
rect 17224 8041 17233 8075
rect 17233 8041 17267 8075
rect 17267 8041 17276 8075
rect 17224 8032 17276 8041
rect 17592 8032 17644 8084
rect 18788 8032 18840 8084
rect 7472 7964 7524 8016
rect 10692 7964 10744 8016
rect 10876 7964 10928 8016
rect 11244 7964 11296 8016
rect 6276 7896 6328 7948
rect 8852 7896 8904 7948
rect 6460 7828 6512 7880
rect 6552 7828 6604 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7104 7828 7156 7880
rect 12256 7896 12308 7948
rect 19064 7964 19116 8016
rect 19524 7964 19576 8016
rect 19984 8075 20036 8084
rect 19984 8041 19993 8075
rect 19993 8041 20027 8075
rect 20027 8041 20036 8075
rect 19984 8032 20036 8041
rect 3976 7760 4028 7812
rect 4068 7803 4120 7812
rect 4068 7769 4077 7803
rect 4077 7769 4111 7803
rect 4111 7769 4120 7803
rect 4068 7760 4120 7769
rect 5356 7760 5408 7812
rect 6368 7692 6420 7744
rect 6460 7692 6512 7744
rect 8024 7760 8076 7812
rect 8484 7803 8536 7812
rect 8484 7769 8493 7803
rect 8493 7769 8527 7803
rect 8527 7769 8536 7803
rect 8484 7760 8536 7769
rect 10784 7760 10836 7812
rect 11428 7828 11480 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 15200 7828 15252 7880
rect 16120 7828 16172 7880
rect 16580 7828 16632 7880
rect 6736 7692 6788 7744
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 10692 7692 10744 7744
rect 11428 7692 11480 7744
rect 12072 7760 12124 7812
rect 13544 7760 13596 7812
rect 14280 7760 14332 7812
rect 15384 7803 15436 7812
rect 15384 7769 15418 7803
rect 15418 7769 15436 7803
rect 15384 7760 15436 7769
rect 17684 7828 17736 7880
rect 19064 7828 19116 7880
rect 18972 7760 19024 7812
rect 16488 7735 16540 7744
rect 16488 7701 16497 7735
rect 16497 7701 16531 7735
rect 16531 7701 16540 7735
rect 16488 7692 16540 7701
rect 19708 7760 19760 7812
rect 19984 7692 20036 7744
rect 7214 7590 7266 7642
rect 7278 7590 7330 7642
rect 7342 7590 7394 7642
rect 7406 7590 7458 7642
rect 7470 7590 7522 7642
rect 13214 7590 13266 7642
rect 13278 7590 13330 7642
rect 13342 7590 13394 7642
rect 13406 7590 13458 7642
rect 13470 7590 13522 7642
rect 19214 7590 19266 7642
rect 19278 7590 19330 7642
rect 19342 7590 19394 7642
rect 19406 7590 19458 7642
rect 19470 7590 19522 7642
rect 4068 7488 4120 7540
rect 2964 7420 3016 7472
rect 5448 7488 5500 7540
rect 5632 7488 5684 7540
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 6552 7488 6604 7540
rect 7104 7420 7156 7472
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 9404 7488 9456 7540
rect 4620 7284 4672 7336
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 5816 7352 5868 7404
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6276 7352 6328 7404
rect 6644 7352 6696 7404
rect 8392 7420 8444 7472
rect 11336 7420 11388 7472
rect 11888 7488 11940 7540
rect 17224 7531 17276 7540
rect 17224 7497 17233 7531
rect 17233 7497 17267 7531
rect 17267 7497 17276 7531
rect 17224 7488 17276 7497
rect 18972 7488 19024 7540
rect 19984 7531 20036 7540
rect 19984 7497 19993 7531
rect 19993 7497 20027 7531
rect 20027 7497 20036 7531
rect 19984 7488 20036 7497
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 7012 7284 7064 7336
rect 6736 7216 6788 7268
rect 7104 7216 7156 7268
rect 7564 7284 7616 7336
rect 2320 7191 2372 7200
rect 2320 7157 2329 7191
rect 2329 7157 2363 7191
rect 2363 7157 2372 7191
rect 2320 7148 2372 7157
rect 3976 7148 4028 7200
rect 5816 7148 5868 7200
rect 7380 7191 7432 7200
rect 7380 7157 7389 7191
rect 7389 7157 7423 7191
rect 7423 7157 7432 7191
rect 7380 7148 7432 7157
rect 10508 7259 10560 7268
rect 10508 7225 10517 7259
rect 10517 7225 10551 7259
rect 10551 7225 10560 7259
rect 10508 7216 10560 7225
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10692 7352 10744 7361
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 10968 7352 11020 7404
rect 15936 7420 15988 7472
rect 16488 7420 16540 7472
rect 19064 7420 19116 7472
rect 11244 7284 11296 7336
rect 12808 7352 12860 7404
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 10876 7216 10928 7268
rect 11796 7216 11848 7268
rect 15476 7148 15528 7200
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 17684 7352 17736 7404
rect 16580 7284 16632 7336
rect 16948 7191 17000 7200
rect 16948 7157 16957 7191
rect 16957 7157 16991 7191
rect 16991 7157 17000 7191
rect 16948 7148 17000 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 10214 7046 10266 7098
rect 10278 7046 10330 7098
rect 10342 7046 10394 7098
rect 10406 7046 10458 7098
rect 10470 7046 10522 7098
rect 16214 7046 16266 7098
rect 16278 7046 16330 7098
rect 16342 7046 16394 7098
rect 16406 7046 16458 7098
rect 16470 7046 16522 7098
rect 5356 6944 5408 6996
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 8392 6944 8444 6996
rect 9864 6944 9916 6996
rect 10968 6944 11020 6996
rect 15200 6944 15252 6996
rect 19064 6944 19116 6996
rect 5448 6808 5500 6860
rect 3976 6740 4028 6792
rect 6092 6740 6144 6792
rect 6460 6740 6512 6792
rect 8024 6808 8076 6860
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7380 6740 7432 6792
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 9772 6808 9824 6860
rect 17040 6876 17092 6928
rect 17316 6851 17368 6860
rect 17316 6817 17325 6851
rect 17325 6817 17359 6851
rect 17359 6817 17368 6851
rect 17316 6808 17368 6817
rect 8484 6740 8536 6792
rect 8852 6740 8904 6792
rect 10876 6740 10928 6792
rect 11152 6783 11204 6792
rect 11152 6749 11161 6783
rect 11161 6749 11195 6783
rect 11195 6749 11204 6783
rect 11152 6740 11204 6749
rect 15476 6783 15528 6792
rect 15476 6749 15510 6783
rect 15510 6749 15528 6783
rect 15476 6740 15528 6749
rect 17684 6740 17736 6792
rect 8392 6672 8444 6724
rect 5540 6604 5592 6656
rect 6736 6604 6788 6656
rect 10784 6672 10836 6724
rect 15568 6672 15620 6724
rect 16580 6647 16632 6656
rect 16580 6613 16589 6647
rect 16589 6613 16623 6647
rect 16623 6613 16632 6647
rect 19616 6672 19668 6724
rect 16580 6604 16632 6613
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 7214 6502 7266 6554
rect 7278 6502 7330 6554
rect 7342 6502 7394 6554
rect 7406 6502 7458 6554
rect 7470 6502 7522 6554
rect 13214 6502 13266 6554
rect 13278 6502 13330 6554
rect 13342 6502 13394 6554
rect 13406 6502 13458 6554
rect 13470 6502 13522 6554
rect 19214 6502 19266 6554
rect 19278 6502 19330 6554
rect 19342 6502 19394 6554
rect 19406 6502 19458 6554
rect 19470 6502 19522 6554
rect 2412 6375 2464 6384
rect 2412 6341 2421 6375
rect 2421 6341 2455 6375
rect 2455 6341 2464 6375
rect 2412 6332 2464 6341
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 1492 6196 1544 6248
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 3056 6239 3108 6248
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 4068 6196 4120 6248
rect 5448 6332 5500 6384
rect 5540 6264 5592 6316
rect 8392 6400 8444 6452
rect 6736 6332 6788 6384
rect 8024 6332 8076 6384
rect 8208 6332 8260 6384
rect 9772 6264 9824 6316
rect 9496 6196 9548 6248
rect 10968 6264 11020 6316
rect 10140 6128 10192 6180
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 2504 6103 2556 6112
rect 2504 6069 2513 6103
rect 2513 6069 2547 6103
rect 2547 6069 2556 6103
rect 2504 6060 2556 6069
rect 4620 6060 4672 6112
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 10784 6060 10836 6112
rect 11520 6060 11572 6112
rect 12164 6196 12216 6248
rect 12348 6307 12400 6316
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 14372 6264 14424 6316
rect 17040 6400 17092 6452
rect 19616 6443 19668 6452
rect 19616 6409 19625 6443
rect 19625 6409 19659 6443
rect 19659 6409 19668 6443
rect 19616 6400 19668 6409
rect 16948 6307 17000 6316
rect 16948 6273 16982 6307
rect 16982 6273 17000 6307
rect 16948 6264 17000 6273
rect 17316 6264 17368 6316
rect 17684 6264 17736 6316
rect 12532 6196 12584 6248
rect 14464 6239 14516 6248
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 14188 6060 14240 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 10214 5958 10266 6010
rect 10278 5958 10330 6010
rect 10342 5958 10394 6010
rect 10406 5958 10458 6010
rect 10470 5958 10522 6010
rect 16214 5958 16266 6010
rect 16278 5958 16330 6010
rect 16342 5958 16394 6010
rect 16406 5958 16458 6010
rect 16470 5958 16522 6010
rect 2044 5856 2096 5908
rect 3056 5856 3108 5908
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 7564 5856 7616 5908
rect 2504 5720 2556 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 3608 5652 3660 5704
rect 4068 5652 4120 5704
rect 8300 5652 8352 5704
rect 8760 5652 8812 5704
rect 9128 5652 9180 5704
rect 9404 5856 9456 5908
rect 10140 5856 10192 5908
rect 10784 5856 10836 5908
rect 12348 5856 12400 5908
rect 14188 5856 14240 5908
rect 17316 5899 17368 5908
rect 17316 5865 17325 5899
rect 17325 5865 17359 5899
rect 17359 5865 17368 5899
rect 17316 5856 17368 5865
rect 13544 5831 13596 5840
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 5908 5627 5960 5636
rect 5908 5593 5917 5627
rect 5917 5593 5951 5627
rect 5951 5593 5960 5627
rect 5908 5584 5960 5593
rect 8024 5584 8076 5636
rect 10876 5652 10928 5704
rect 9680 5584 9732 5636
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 8392 5516 8444 5568
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 9404 5516 9456 5568
rect 13544 5652 13596 5704
rect 15108 5720 15160 5772
rect 15844 5695 15896 5704
rect 15844 5661 15853 5695
rect 15853 5661 15887 5695
rect 15887 5661 15896 5695
rect 15844 5652 15896 5661
rect 16580 5652 16632 5704
rect 11152 5516 11204 5568
rect 11520 5516 11572 5568
rect 12624 5559 12676 5568
rect 12624 5525 12633 5559
rect 12633 5525 12667 5559
rect 12667 5525 12676 5559
rect 12624 5516 12676 5525
rect 7214 5414 7266 5466
rect 7278 5414 7330 5466
rect 7342 5414 7394 5466
rect 7406 5414 7458 5466
rect 7470 5414 7522 5466
rect 13214 5414 13266 5466
rect 13278 5414 13330 5466
rect 13342 5414 13394 5466
rect 13406 5414 13458 5466
rect 13470 5414 13522 5466
rect 19214 5414 19266 5466
rect 19278 5414 19330 5466
rect 19342 5414 19394 5466
rect 19406 5414 19458 5466
rect 19470 5414 19522 5466
rect 2044 5312 2096 5364
rect 2688 5312 2740 5364
rect 2780 5312 2832 5364
rect 4804 5312 4856 5364
rect 1400 5176 1452 5228
rect 2320 5287 2372 5296
rect 2320 5253 2329 5287
rect 2329 5253 2363 5287
rect 2363 5253 2372 5287
rect 2320 5244 2372 5253
rect 3148 5108 3200 5160
rect 1584 5040 1636 5092
rect 4620 5244 4672 5296
rect 3700 5108 3752 5160
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 7104 5312 7156 5364
rect 8668 5312 8720 5364
rect 9680 5312 9732 5364
rect 12808 5355 12860 5364
rect 12808 5321 12817 5355
rect 12817 5321 12851 5355
rect 12851 5321 12860 5355
rect 12808 5312 12860 5321
rect 14372 5312 14424 5364
rect 14464 5312 14516 5364
rect 8300 5244 8352 5296
rect 3424 5040 3476 5092
rect 4068 5040 4120 5092
rect 8208 5176 8260 5228
rect 9312 5244 9364 5296
rect 11152 5244 11204 5296
rect 11336 5244 11388 5296
rect 13912 5244 13964 5296
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 8852 5219 8904 5228
rect 8852 5185 8889 5219
rect 8889 5185 8904 5219
rect 8852 5176 8904 5185
rect 3332 5015 3384 5024
rect 3332 4981 3341 5015
rect 3341 4981 3375 5015
rect 3375 4981 3384 5015
rect 3332 4972 3384 4981
rect 6460 5151 6512 5160
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6460 5108 6512 5117
rect 9404 5176 9456 5228
rect 11244 5219 11296 5228
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 4712 4972 4764 5024
rect 8208 5015 8260 5024
rect 8208 4981 8217 5015
rect 8217 4981 8251 5015
rect 8251 4981 8260 5015
rect 8208 4972 8260 4981
rect 12532 5108 12584 5160
rect 20812 5176 20864 5228
rect 13268 5040 13320 5092
rect 11060 5015 11112 5024
rect 11060 4981 11069 5015
rect 11069 4981 11103 5015
rect 11103 4981 11112 5015
rect 11060 4972 11112 4981
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 10214 4870 10266 4922
rect 10278 4870 10330 4922
rect 10342 4870 10394 4922
rect 10406 4870 10458 4922
rect 10470 4870 10522 4922
rect 16214 4870 16266 4922
rect 16278 4870 16330 4922
rect 16342 4870 16394 4922
rect 16406 4870 16458 4922
rect 16470 4870 16522 4922
rect 4712 4768 4764 4820
rect 4804 4768 4856 4820
rect 5908 4768 5960 4820
rect 6460 4768 6512 4820
rect 11704 4768 11756 4820
rect 3700 4564 3752 4616
rect 3792 4496 3844 4548
rect 4160 4564 4212 4616
rect 4620 4564 4672 4616
rect 9128 4700 9180 4752
rect 13268 4768 13320 4820
rect 13360 4768 13412 4820
rect 8300 4564 8352 4616
rect 8392 4564 8444 4616
rect 8484 4496 8536 4548
rect 9220 4496 9272 4548
rect 10876 4539 10928 4548
rect 10876 4505 10885 4539
rect 10885 4505 10919 4539
rect 10919 4505 10928 4539
rect 12624 4564 12676 4616
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 10876 4496 10928 4505
rect 8392 4428 8444 4480
rect 8760 4428 8812 4480
rect 9772 4428 9824 4480
rect 12900 4428 12952 4480
rect 13544 4428 13596 4480
rect 13728 4471 13780 4480
rect 13728 4437 13737 4471
rect 13737 4437 13771 4471
rect 13771 4437 13780 4471
rect 13728 4428 13780 4437
rect 7214 4326 7266 4378
rect 7278 4326 7330 4378
rect 7342 4326 7394 4378
rect 7406 4326 7458 4378
rect 7470 4326 7522 4378
rect 13214 4326 13266 4378
rect 13278 4326 13330 4378
rect 13342 4326 13394 4378
rect 13406 4326 13458 4378
rect 13470 4326 13522 4378
rect 19214 4326 19266 4378
rect 19278 4326 19330 4378
rect 19342 4326 19394 4378
rect 19406 4326 19458 4378
rect 19470 4326 19522 4378
rect 9128 4224 9180 4276
rect 12532 4224 12584 4276
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8392 4088 8444 4140
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 3792 3952 3844 4004
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 7012 3884 7064 3936
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 8852 4088 8904 4140
rect 9128 4088 9180 4140
rect 9220 4131 9272 4140
rect 9220 4097 9229 4131
rect 9229 4097 9263 4131
rect 9263 4097 9272 4131
rect 9220 4088 9272 4097
rect 9588 4088 9640 4140
rect 11060 4156 11112 4208
rect 13728 4224 13780 4276
rect 14372 4156 14424 4208
rect 10968 4088 11020 4140
rect 12900 4088 12952 4140
rect 9220 3952 9272 4004
rect 9496 3952 9548 4004
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 9680 3884 9732 3936
rect 12808 3884 12860 3936
rect 14832 3927 14884 3936
rect 14832 3893 14841 3927
rect 14841 3893 14875 3927
rect 14875 3893 14884 3927
rect 14832 3884 14884 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 10214 3782 10266 3834
rect 10278 3782 10330 3834
rect 10342 3782 10394 3834
rect 10406 3782 10458 3834
rect 10470 3782 10522 3834
rect 16214 3782 16266 3834
rect 16278 3782 16330 3834
rect 16342 3782 16394 3834
rect 16406 3782 16458 3834
rect 16470 3782 16522 3834
rect 20 3680 72 3732
rect 1400 3680 1452 3732
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 4068 3680 4120 3732
rect 8852 3680 8904 3732
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 12440 3680 12492 3732
rect 8024 3544 8076 3596
rect 8300 3544 8352 3596
rect 3608 3476 3660 3528
rect 4344 3476 4396 3528
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 8576 3476 8628 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9220 3476 9272 3528
rect 9588 3519 9640 3528
rect 9588 3485 9591 3519
rect 9591 3485 9640 3519
rect 9588 3476 9640 3485
rect 5448 3451 5500 3460
rect 5448 3417 5457 3451
rect 5457 3417 5491 3451
rect 5491 3417 5500 3451
rect 5448 3408 5500 3417
rect 8944 3340 8996 3392
rect 9312 3451 9364 3460
rect 9312 3417 9321 3451
rect 9321 3417 9355 3451
rect 9355 3417 9364 3451
rect 9312 3408 9364 3417
rect 11520 3408 11572 3460
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 9956 3383 10008 3392
rect 9956 3349 9965 3383
rect 9965 3349 9999 3383
rect 9999 3349 10008 3383
rect 9956 3340 10008 3349
rect 12532 3408 12584 3460
rect 13820 3680 13872 3732
rect 14740 3680 14792 3732
rect 13544 3655 13596 3664
rect 13544 3621 13553 3655
rect 13553 3621 13587 3655
rect 13587 3621 13596 3655
rect 13544 3612 13596 3621
rect 14832 3544 14884 3596
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 11796 3383 11848 3392
rect 11796 3349 11805 3383
rect 11805 3349 11839 3383
rect 11839 3349 11848 3383
rect 11796 3340 11848 3349
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 14372 3408 14424 3460
rect 14832 3408 14884 3460
rect 7214 3238 7266 3290
rect 7278 3238 7330 3290
rect 7342 3238 7394 3290
rect 7406 3238 7458 3290
rect 7470 3238 7522 3290
rect 13214 3238 13266 3290
rect 13278 3238 13330 3290
rect 13342 3238 13394 3290
rect 13406 3238 13458 3290
rect 13470 3238 13522 3290
rect 19214 3238 19266 3290
rect 19278 3238 19330 3290
rect 19342 3238 19394 3290
rect 19406 3238 19458 3290
rect 19470 3238 19522 3290
rect 5448 3136 5500 3188
rect 8392 3136 8444 3188
rect 9220 3136 9272 3188
rect 9956 3136 10008 3188
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 12716 3136 12768 3188
rect 3332 3068 3384 3120
rect 4344 3068 4396 3120
rect 9404 3068 9456 3120
rect 13728 3136 13780 3188
rect 14740 3136 14792 3188
rect 8944 3000 8996 3052
rect 14280 3068 14332 3120
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12440 3000 12492 3009
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 10416 2975 10468 2984
rect 10416 2941 10425 2975
rect 10425 2941 10459 2975
rect 10459 2941 10468 2975
rect 10416 2932 10468 2941
rect 3792 2796 3844 2848
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 14372 2975 14424 2984
rect 14372 2941 14381 2975
rect 14381 2941 14415 2975
rect 14415 2941 14424 2975
rect 14372 2932 14424 2941
rect 20628 2864 20680 2916
rect 12348 2839 12400 2848
rect 12348 2805 12357 2839
rect 12357 2805 12391 2839
rect 12391 2805 12400 2839
rect 12348 2796 12400 2805
rect 13544 2796 13596 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 10214 2694 10266 2746
rect 10278 2694 10330 2746
rect 10342 2694 10394 2746
rect 10406 2694 10458 2746
rect 10470 2694 10522 2746
rect 16214 2694 16266 2746
rect 16278 2694 16330 2746
rect 16342 2694 16394 2746
rect 16406 2694 16458 2746
rect 16470 2694 16522 2746
rect 10968 2592 11020 2644
rect 11244 2592 11296 2644
rect 12072 2592 12124 2644
rect 12532 2592 12584 2644
rect 14372 2592 14424 2644
rect 10048 2524 10100 2576
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 12348 2456 12400 2508
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 9772 2388 9824 2440
rect 10876 2388 10928 2440
rect 11796 2388 11848 2440
rect 12256 2388 12308 2440
rect 12440 2388 12492 2440
rect 14096 2524 14148 2576
rect 15200 2388 15252 2440
rect 15568 2363 15620 2372
rect 15568 2329 15577 2363
rect 15577 2329 15611 2363
rect 15611 2329 15620 2363
rect 15568 2320 15620 2329
rect 7214 2150 7266 2202
rect 7278 2150 7330 2202
rect 7342 2150 7394 2202
rect 7406 2150 7458 2202
rect 7470 2150 7522 2202
rect 13214 2150 13266 2202
rect 13278 2150 13330 2202
rect 13342 2150 13394 2202
rect 13406 2150 13458 2202
rect 13470 2150 13522 2202
rect 19214 2150 19266 2202
rect 19278 2150 19330 2202
rect 19342 2150 19394 2202
rect 19406 2150 19458 2202
rect 19470 2150 19522 2202
<< metal2 >>
rect 3238 23290 3294 24090
rect 8390 23290 8446 24090
rect 13542 23290 13598 24090
rect 18694 23290 18750 24090
rect 3252 21554 3280 23290
rect 3606 21856 3662 21865
rect 3606 21791 3662 21800
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3528 19378 3556 19654
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 2792 18766 2820 19314
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 2056 18426 2084 18566
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1400 17536 1452 17542
rect 1400 17478 1452 17484
rect 1412 17202 1440 17478
rect 1688 17338 1716 17614
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 952 16425 980 16458
rect 938 16416 994 16425
rect 938 16351 994 16360
rect 1412 16114 1440 17138
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 12782 1440 16050
rect 1688 16046 1716 16390
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1688 15502 1716 15982
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 15162 1716 15438
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1688 14618 1716 14894
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1780 14414 1808 14758
rect 1872 14414 1900 15302
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1596 13802 1624 14350
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12238 1440 12718
rect 1676 12708 1728 12714
rect 1676 12650 1728 12656
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11762 1440 12174
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1596 11898 1624 12038
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1688 11354 1716 12650
rect 1768 12640 1820 12646
rect 1768 12582 1820 12588
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1780 12434 1808 12582
rect 1964 12442 1992 12582
rect 1952 12436 2004 12442
rect 1780 12406 1900 12434
rect 1872 12238 1900 12406
rect 1952 12378 2004 12384
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 9586 1624 10406
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 9178 1808 9318
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1780 7886 1808 8230
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1504 5386 1532 6190
rect 2056 5914 2084 16594
rect 2148 12434 2176 18022
rect 2688 17604 2740 17610
rect 2688 17546 2740 17552
rect 2700 17338 2728 17546
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 2688 16516 2740 16522
rect 2688 16458 2740 16464
rect 2700 16250 2728 16458
rect 3528 16454 3556 16934
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 3344 16114 3372 16390
rect 3436 16182 3464 16390
rect 3528 16182 3556 16390
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3516 16176 3568 16182
rect 3516 16118 3568 16124
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3528 15638 3556 16118
rect 3516 15632 3568 15638
rect 3516 15574 3568 15580
rect 3528 15094 3556 15574
rect 3516 15088 3568 15094
rect 3516 15030 3568 15036
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3160 14618 3188 14758
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3344 14074 3372 14962
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3528 14006 3556 14758
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2700 13326 2728 13738
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2516 12850 2544 13126
rect 2700 12986 2728 13262
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12986 3188 13126
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2516 12434 2544 12786
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 2148 12406 2268 12434
rect 2516 12406 2636 12434
rect 2240 10674 2268 12406
rect 2608 12306 2636 12406
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 3240 12232 3292 12238
rect 3436 12220 3464 12718
rect 3528 12442 3556 13262
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3292 12192 3464 12220
rect 3240 12174 3292 12180
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2424 11898 2452 12106
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 3436 11762 3464 12192
rect 3528 12170 3556 12378
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 3436 9994 3464 11698
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9722 2820 9862
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8634 2268 8774
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1412 5358 1532 5386
rect 1412 5234 1440 5358
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 3738 1440 5170
rect 1596 5098 1624 5510
rect 2056 5370 2084 5850
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2332 5302 2360 7142
rect 2516 6914 2544 7754
rect 2976 7478 3004 8230
rect 3620 8090 3648 21791
rect 7214 21788 7522 21797
rect 7214 21786 7220 21788
rect 7276 21786 7300 21788
rect 7356 21786 7380 21788
rect 7436 21786 7460 21788
rect 7516 21786 7522 21788
rect 7276 21734 7278 21786
rect 7458 21734 7460 21786
rect 7214 21732 7220 21734
rect 7276 21732 7300 21734
rect 7356 21732 7380 21734
rect 7436 21732 7460 21734
rect 7516 21732 7522 21734
rect 7214 21723 7522 21732
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4540 20466 4568 20742
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 20058 3924 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 5000 18970 5028 19314
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 3804 15978 3832 17614
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4264 17134 4292 17478
rect 4632 17338 4660 17478
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4344 17128 4396 17134
rect 4816 17116 4844 17614
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 4396 17088 4844 17116
rect 4344 17070 4396 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3896 16046 3924 16730
rect 4632 16454 4660 17088
rect 5092 16522 5120 17478
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16590 5304 16934
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4908 16114 4936 16390
rect 5092 16114 5120 16458
rect 5276 16250 5304 16526
rect 5368 16250 5396 17614
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5552 16522 5580 17478
rect 5644 17202 5672 17478
rect 5736 17202 5764 21422
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6288 20398 6316 20946
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6288 20058 6316 20334
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6092 19712 6144 19718
rect 6092 19654 6144 19660
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6104 18834 6132 19654
rect 6196 19242 6224 19654
rect 6288 19514 6316 19994
rect 6932 19854 6960 21490
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7300 21010 7328 21286
rect 7576 21010 7604 21286
rect 7668 21146 7696 21286
rect 8404 21146 8432 23290
rect 13556 22094 13584 23290
rect 13556 22066 13860 22094
rect 13214 21788 13522 21797
rect 13214 21786 13220 21788
rect 13276 21786 13300 21788
rect 13356 21786 13380 21788
rect 13436 21786 13460 21788
rect 13516 21786 13522 21788
rect 13276 21734 13278 21786
rect 13458 21734 13460 21786
rect 13214 21732 13220 21734
rect 13276 21732 13300 21734
rect 13356 21732 13380 21734
rect 13436 21732 13460 21734
rect 13516 21732 13522 21734
rect 13214 21723 13522 21732
rect 13832 21622 13860 22066
rect 13820 21616 13872 21622
rect 13820 21558 13872 21564
rect 18708 21554 18736 23290
rect 19214 21788 19522 21797
rect 19214 21786 19220 21788
rect 19276 21786 19300 21788
rect 19356 21786 19380 21788
rect 19436 21786 19460 21788
rect 19516 21786 19522 21788
rect 19276 21734 19278 21786
rect 19458 21734 19460 21786
rect 19214 21732 19220 21734
rect 19276 21732 19300 21734
rect 19356 21732 19380 21734
rect 19436 21732 19460 21734
rect 19516 21732 19522 21734
rect 19214 21723 19522 21732
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10060 21146 10088 21422
rect 10214 21244 10522 21253
rect 10214 21242 10220 21244
rect 10276 21242 10300 21244
rect 10356 21242 10380 21244
rect 10436 21242 10460 21244
rect 10516 21242 10522 21244
rect 10276 21190 10278 21242
rect 10458 21190 10460 21242
rect 10214 21188 10220 21190
rect 10276 21188 10300 21190
rect 10356 21188 10380 21190
rect 10436 21188 10460 21190
rect 10516 21188 10522 21190
rect 10214 21179 10522 21188
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7564 21004 7616 21010
rect 7564 20946 7616 20952
rect 10888 20942 10916 21422
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 7214 20700 7522 20709
rect 7214 20698 7220 20700
rect 7276 20698 7300 20700
rect 7356 20698 7380 20700
rect 7436 20698 7460 20700
rect 7516 20698 7522 20700
rect 7276 20646 7278 20698
rect 7458 20646 7460 20698
rect 7214 20644 7220 20646
rect 7276 20644 7300 20646
rect 7356 20644 7380 20646
rect 7436 20644 7460 20646
rect 7516 20644 7522 20646
rect 7214 20635 7522 20644
rect 8496 20602 8524 20742
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6380 19514 6408 19722
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6184 19236 6236 19242
rect 6184 19178 6236 19184
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6104 17746 6132 18770
rect 6196 18766 6224 19178
rect 6380 18970 6408 19450
rect 6932 18970 6960 19790
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 7024 18834 7052 20198
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7214 19612 7522 19621
rect 7214 19610 7220 19612
rect 7276 19610 7300 19612
rect 7356 19610 7380 19612
rect 7436 19610 7460 19612
rect 7516 19610 7522 19612
rect 7276 19558 7278 19610
rect 7458 19558 7460 19610
rect 7214 19556 7220 19558
rect 7276 19556 7300 19558
rect 7356 19556 7380 19558
rect 7436 19556 7460 19558
rect 7516 19556 7522 19558
rect 7214 19547 7522 19556
rect 7576 19446 7604 19654
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7852 18834 7880 19246
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 7024 18426 7052 18770
rect 8312 18766 8340 20470
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8404 20058 8432 20334
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8588 19854 8616 20198
rect 9416 19922 9444 20742
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8588 19514 8616 19790
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8588 18698 8616 19450
rect 9600 19378 9628 20878
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 20262 9720 20742
rect 11532 20534 11560 21490
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8772 18970 8800 19178
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 8576 18692 8628 18698
rect 8576 18634 8628 18640
rect 7214 18524 7522 18533
rect 7214 18522 7220 18524
rect 7276 18522 7300 18524
rect 7356 18522 7380 18524
rect 7436 18522 7460 18524
rect 7516 18522 7522 18524
rect 7276 18470 7278 18522
rect 7458 18470 7460 18522
rect 7214 18468 7220 18470
rect 7276 18468 7300 18470
rect 7356 18468 7380 18470
rect 7436 18468 7460 18470
rect 7516 18468 7522 18470
rect 7214 18459 7522 18468
rect 7576 18426 7604 18634
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 7214 17436 7522 17445
rect 7214 17434 7220 17436
rect 7276 17434 7300 17436
rect 7356 17434 7380 17436
rect 7436 17434 7460 17436
rect 7516 17434 7522 17436
rect 7276 17382 7278 17434
rect 7458 17382 7460 17434
rect 7214 17380 7220 17382
rect 7276 17380 7300 17382
rect 7356 17380 7380 17382
rect 7436 17380 7460 17382
rect 7516 17380 7522 17382
rect 7214 17371 7522 17380
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6196 16794 6224 16934
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6656 16522 6684 17138
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6840 16454 6868 17138
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7668 16794 7696 17070
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 5080 16108 5132 16114
rect 5080 16050 5132 16056
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3792 15972 3844 15978
rect 3792 15914 3844 15920
rect 3896 15094 3924 15982
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 6092 15632 6144 15638
rect 6092 15574 6144 15580
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3884 15088 3936 15094
rect 3884 15030 3936 15036
rect 3804 13938 3832 15030
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 3988 14618 4016 14962
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3988 14074 4016 14554
rect 4080 14346 4108 14962
rect 6012 14958 6040 15302
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 4080 13870 4108 14282
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3976 12844 4028 12850
rect 4080 12832 4108 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4028 12804 4108 12832
rect 3976 12786 4028 12792
rect 4172 12730 4200 13126
rect 4356 12986 4384 13126
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4540 12866 4568 13330
rect 4540 12838 4660 12866
rect 4080 12702 4200 12730
rect 4080 12170 4108 12702
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4080 11898 4108 12106
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 10810 4660 12838
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12238 4752 12582
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4816 10674 4844 10746
rect 5184 10742 5212 14282
rect 5736 14074 5764 14894
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5828 14074 5856 14350
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 6104 13938 6132 15574
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14074 6408 14758
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5368 12442 5396 13806
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5460 12782 5488 13330
rect 5644 12832 5672 13874
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13530 6040 13670
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6380 12986 6408 13262
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 5724 12844 5776 12850
rect 5644 12804 5724 12832
rect 5724 12786 5776 12792
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 5276 11354 5304 12106
rect 6840 11694 6868 16390
rect 7214 16348 7522 16357
rect 7214 16346 7220 16348
rect 7276 16346 7300 16348
rect 7356 16346 7380 16348
rect 7436 16346 7460 16348
rect 7516 16346 7522 16348
rect 7276 16294 7278 16346
rect 7458 16294 7460 16346
rect 7214 16292 7220 16294
rect 7276 16292 7300 16294
rect 7356 16292 7380 16294
rect 7436 16292 7460 16294
rect 7516 16292 7522 16294
rect 7214 16283 7522 16292
rect 8312 15910 8340 16390
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 7024 15162 7052 15302
rect 7214 15260 7522 15269
rect 7214 15258 7220 15260
rect 7276 15258 7300 15260
rect 7356 15258 7380 15260
rect 7436 15258 7460 15260
rect 7516 15258 7522 15260
rect 7276 15206 7278 15258
rect 7458 15206 7460 15258
rect 7214 15204 7220 15206
rect 7276 15204 7300 15206
rect 7356 15204 7380 15206
rect 7436 15204 7460 15206
rect 7516 15204 7522 15206
rect 7214 15195 7522 15204
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7668 14482 7696 14758
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7760 14346 7788 14962
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 6932 14006 6960 14282
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7214 14172 7522 14181
rect 7214 14170 7220 14172
rect 7276 14170 7300 14172
rect 7356 14170 7380 14172
rect 7436 14170 7460 14172
rect 7516 14170 7522 14172
rect 7276 14118 7278 14170
rect 7458 14118 7460 14170
rect 7214 14116 7220 14118
rect 7276 14116 7300 14118
rect 7356 14116 7380 14118
rect 7436 14116 7460 14118
rect 7516 14116 7522 14118
rect 7214 14107 7522 14116
rect 7668 14074 7696 14214
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 7760 13326 7788 14282
rect 7852 14006 7880 15370
rect 7944 14482 7972 15846
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7852 13530 7880 13942
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5276 11218 5304 11290
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 6932 11150 6960 13126
rect 7214 13084 7522 13093
rect 7214 13082 7220 13084
rect 7276 13082 7300 13084
rect 7356 13082 7380 13084
rect 7436 13082 7460 13084
rect 7516 13082 7522 13084
rect 7276 13030 7278 13082
rect 7458 13030 7460 13082
rect 7214 13028 7220 13030
rect 7276 13028 7300 13030
rect 7356 13028 7380 13030
rect 7436 13028 7460 13030
rect 7516 13028 7522 13030
rect 7214 13019 7522 13028
rect 7944 12986 7972 14418
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10810 5580 11018
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 7024 10674 7052 10950
rect 7116 10810 7144 12854
rect 7214 11996 7522 12005
rect 7214 11994 7220 11996
rect 7276 11994 7300 11996
rect 7356 11994 7380 11996
rect 7436 11994 7460 11996
rect 7516 11994 7522 11996
rect 7276 11942 7278 11994
rect 7458 11942 7460 11994
rect 7214 11940 7220 11942
rect 7276 11940 7300 11942
rect 7356 11940 7380 11942
rect 7436 11940 7460 11942
rect 7516 11940 7522 11942
rect 7214 11931 7522 11940
rect 7944 11354 7972 12922
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7214 10908 7522 10917
rect 7214 10906 7220 10908
rect 7276 10906 7300 10908
rect 7356 10906 7380 10908
rect 7436 10906 7460 10908
rect 7516 10906 7522 10908
rect 7276 10854 7278 10906
rect 7458 10854 7460 10906
rect 7214 10852 7220 10854
rect 7276 10852 7300 10854
rect 7356 10852 7380 10854
rect 7436 10852 7460 10854
rect 7516 10852 7522 10854
rect 7214 10843 7522 10852
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 5540 10668 5592 10674
rect 7012 10668 7064 10674
rect 5540 10610 5592 10616
rect 6932 10628 7012 10656
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4816 10266 4844 10610
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 3988 9382 4016 9930
rect 4356 9722 4384 9930
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4816 9450 4844 10202
rect 4908 9722 4936 10542
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5092 9722 5120 10406
rect 5552 10266 5580 10610
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3988 7818 4016 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9024 4660 9318
rect 4448 8996 4660 9024
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4264 8566 4292 8774
rect 4448 8566 4476 8996
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4632 8430 4660 8842
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4724 8566 4752 8774
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 3988 7206 4016 7754
rect 4080 7546 4108 7754
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4632 7342 4660 8366
rect 4908 8294 4936 9522
rect 5092 9382 5120 9522
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5184 8498 5212 8910
rect 5368 8906 5396 9386
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5460 8838 5488 9318
rect 5552 9178 5580 10202
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 5644 9722 5672 9862
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 6656 9586 6684 9862
rect 6748 9586 6776 10542
rect 6932 10146 6960 10628
rect 7012 10610 7064 10616
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6840 10118 6960 10146
rect 6840 9722 6868 10118
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6932 9722 6960 9930
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5644 9042 5672 9318
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5276 8634 5304 8774
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7410 5212 8230
rect 5276 7410 5304 8570
rect 5644 8498 5672 8978
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5644 8362 5672 8434
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 2424 6886 2544 6914
rect 2424 6390 2452 6886
rect 3988 6798 4016 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5368 7002 5396 7754
rect 5460 7546 5488 7822
rect 5644 7546 5672 7958
rect 5736 7546 5764 9454
rect 5828 9178 5856 9454
rect 5920 9178 5948 9522
rect 6656 9450 6684 9522
rect 6748 9450 6776 9522
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 7024 9178 7052 10202
rect 7116 9654 7144 10406
rect 7484 10130 7512 10610
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7214 9820 7522 9829
rect 7214 9818 7220 9820
rect 7276 9818 7300 9820
rect 7356 9818 7380 9820
rect 7436 9818 7460 9820
rect 7516 9818 7522 9820
rect 7276 9766 7278 9818
rect 7458 9766 7460 9818
rect 7214 9764 7220 9766
rect 7276 9764 7300 9766
rect 7356 9764 7380 9766
rect 7436 9764 7460 9766
rect 7516 9764 7522 9766
rect 7214 9755 7522 9764
rect 7576 9722 7604 10474
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7104 9648 7156 9654
rect 7668 9602 7696 10746
rect 7944 10606 7972 11290
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7760 10266 7788 10542
rect 8036 10266 8064 10610
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7104 9590 7156 9596
rect 7576 9574 7696 9602
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7116 9178 7144 9454
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 5828 8634 5856 9114
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5828 8090 5856 8434
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5460 6866 5488 7482
rect 5828 7410 5856 8026
rect 5920 7410 5948 8434
rect 6288 8362 6316 8910
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6276 8356 6328 8362
rect 6276 8298 6328 8304
rect 6288 7954 6316 8298
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6380 7750 6408 8230
rect 6472 8022 6500 8774
rect 7024 8634 7052 9114
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6656 8294 6684 8434
rect 6932 8378 6960 8502
rect 6736 8356 6788 8362
rect 6932 8350 7052 8378
rect 6736 8298 6788 8304
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6472 7886 6500 7958
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 5828 7206 5856 7346
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 5460 6390 5488 6802
rect 6104 6798 6132 7278
rect 6288 7002 6316 7346
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6472 6798 6500 7686
rect 6564 7546 6592 7822
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6656 7410 6684 8230
rect 6748 7886 6776 8298
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 7024 7750 7052 8350
rect 7116 7886 7144 9114
rect 7576 8906 7604 9574
rect 7760 9178 7788 10066
rect 8036 9926 8064 10202
rect 8128 10062 8156 10950
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7944 9450 7972 9522
rect 8220 9518 8248 11018
rect 8208 9512 8260 9518
rect 8128 9460 8208 9466
rect 8128 9454 8260 9460
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 8128 9438 8248 9454
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7214 8732 7522 8741
rect 7214 8730 7220 8732
rect 7276 8730 7300 8732
rect 7356 8730 7380 8732
rect 7436 8730 7460 8732
rect 7516 8730 7522 8732
rect 7276 8678 7278 8730
rect 7458 8678 7460 8730
rect 7214 8676 7220 8678
rect 7276 8676 7300 8678
rect 7356 8676 7380 8678
rect 7436 8676 7460 8678
rect 7516 8676 7522 8678
rect 7214 8667 7522 8676
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7484 8022 7512 8230
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6748 7274 6776 7686
rect 7024 7342 7052 7686
rect 7116 7478 7144 7822
rect 7214 7644 7522 7653
rect 7214 7642 7220 7644
rect 7276 7642 7300 7644
rect 7356 7642 7380 7644
rect 7436 7642 7460 7644
rect 7516 7642 7522 7644
rect 7276 7590 7278 7642
rect 7458 7590 7460 7642
rect 7214 7588 7220 7590
rect 7276 7588 7300 7590
rect 7356 7588 7380 7590
rect 7436 7588 7460 7590
rect 7516 7588 7522 7590
rect 7214 7579 7522 7588
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7576 7342 7604 8842
rect 7852 8838 7880 9318
rect 7944 8974 7972 9386
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 7818 8064 8774
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 6748 6798 6776 7210
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5552 6322 5580 6598
rect 6748 6390 6776 6598
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2516 5778 2544 6054
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2700 5370 2728 6258
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 2792 5370 2820 6190
rect 3068 5914 3096 6190
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 4080 5710 4108 6190
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 3148 5160 3200 5166
rect 3200 5108 3464 5114
rect 3148 5102 3464 5108
rect 3160 5098 3464 5102
rect 1584 5092 1636 5098
rect 3160 5092 3476 5098
rect 3160 5086 3424 5092
rect 1584 5034 1636 5040
rect 3424 5034 3476 5040
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 20 3732 72 3738
rect 20 3674 72 3680
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 32 800 60 3674
rect 3344 3126 3372 4966
rect 3620 3534 3648 5646
rect 4632 5302 4660 6054
rect 5552 5914 5580 6258
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5908 5636 5960 5642
rect 5908 5578 5960 5584
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4620 5296 4672 5302
rect 3896 5234 4108 5250
rect 4620 5238 4672 5244
rect 3896 5228 4120 5234
rect 3896 5222 4068 5228
rect 3700 5160 3752 5166
rect 3896 5114 3924 5222
rect 4068 5170 4120 5176
rect 3700 5102 3752 5108
rect 3712 4622 3740 5102
rect 3804 5086 3924 5114
rect 4068 5092 4120 5098
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3804 4554 3832 5086
rect 4068 5034 4120 5040
rect 4080 4604 4108 5034
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4622 4660 5238
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4826 4752 4966
rect 4816 4826 4844 5306
rect 5920 4826 5948 5578
rect 7116 5370 7144 7210
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 6798 7420 7142
rect 8036 6866 8064 7754
rect 8128 7546 8156 9438
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8566 8248 8910
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7214 6556 7522 6565
rect 7214 6554 7220 6556
rect 7276 6554 7300 6556
rect 7356 6554 7380 6556
rect 7436 6554 7460 6556
rect 7516 6554 7522 6556
rect 7276 6502 7278 6554
rect 7458 6502 7460 6554
rect 7214 6500 7220 6502
rect 7276 6500 7300 6502
rect 7356 6500 7380 6502
rect 7436 6500 7460 6502
rect 7516 6500 7522 6502
rect 7214 6491 7522 6500
rect 7576 5914 7604 6734
rect 8036 6390 8064 6802
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6390 8248 6734
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 8036 5642 8064 6326
rect 8312 5710 8340 13670
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8404 12442 8432 12718
rect 8392 12436 8444 12442
rect 8588 12434 8616 16934
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8680 16454 8708 16526
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8864 16182 8892 18770
rect 9048 18426 9076 19110
rect 9140 18970 9168 19314
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9220 19236 9272 19242
rect 9220 19178 9272 19184
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9128 18692 9180 18698
rect 9128 18634 9180 18640
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9140 18358 9168 18634
rect 9232 18426 9260 19178
rect 9324 18766 9352 19246
rect 9600 18970 9628 19314
rect 9692 19310 9720 20198
rect 10060 20058 10088 20334
rect 10214 20156 10522 20165
rect 10214 20154 10220 20156
rect 10276 20154 10300 20156
rect 10356 20154 10380 20156
rect 10436 20154 10460 20156
rect 10516 20154 10522 20156
rect 10276 20102 10278 20154
rect 10458 20102 10460 20154
rect 10214 20100 10220 20102
rect 10276 20100 10300 20102
rect 10356 20100 10380 20102
rect 10436 20100 10460 20102
rect 10516 20100 10522 20102
rect 10214 20091 10522 20100
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 11532 19854 11560 20470
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11532 19514 11560 19790
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9496 18896 9548 18902
rect 9496 18838 9548 18844
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9128 18352 9180 18358
rect 9128 18294 9180 18300
rect 9324 18086 9352 18702
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9416 18426 9444 18566
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9508 18290 9536 18838
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9600 18222 9628 18906
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9784 18426 9812 18634
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 10060 18290 10088 19110
rect 10214 19068 10522 19077
rect 10214 19066 10220 19068
rect 10276 19066 10300 19068
rect 10356 19066 10380 19068
rect 10436 19066 10460 19068
rect 10516 19066 10522 19068
rect 10276 19014 10278 19066
rect 10458 19014 10460 19066
rect 10214 19012 10220 19014
rect 10276 19012 10300 19014
rect 10356 19012 10380 19014
rect 10436 19012 10460 19014
rect 10516 19012 10522 19014
rect 10214 19003 10522 19012
rect 11164 18970 11192 19246
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11532 18834 11560 19450
rect 12360 19446 12388 20198
rect 12452 19854 12480 20742
rect 13214 20700 13522 20709
rect 13214 20698 13220 20700
rect 13276 20698 13300 20700
rect 13356 20698 13380 20700
rect 13436 20698 13460 20700
rect 13516 20698 13522 20700
rect 13276 20646 13278 20698
rect 13458 20646 13460 20698
rect 13214 20644 13220 20646
rect 13276 20644 13300 20646
rect 13356 20644 13380 20646
rect 13436 20644 13460 20646
rect 13516 20644 13522 20646
rect 13214 20635 13522 20644
rect 13832 20534 13860 20878
rect 14292 20806 14320 21286
rect 16214 21244 16522 21253
rect 16214 21242 16220 21244
rect 16276 21242 16300 21244
rect 16356 21242 16380 21244
rect 16436 21242 16460 21244
rect 16516 21242 16522 21244
rect 16276 21190 16278 21242
rect 16458 21190 16460 21242
rect 16214 21188 16220 21190
rect 16276 21188 16300 21190
rect 16356 21188 16380 21190
rect 16436 21188 16460 21190
rect 16516 21188 16522 21190
rect 16214 21179 16522 21188
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13464 20058 13492 20402
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 13464 19802 13492 19994
rect 13636 19848 13688 19854
rect 13464 19774 13584 19802
rect 13636 19790 13688 19796
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 13214 19612 13522 19621
rect 13214 19610 13220 19612
rect 13276 19610 13300 19612
rect 13356 19610 13380 19612
rect 13436 19610 13460 19612
rect 13516 19610 13522 19612
rect 13276 19558 13278 19610
rect 13458 19558 13460 19610
rect 13214 19556 13220 19558
rect 13276 19556 13300 19558
rect 13356 19556 13380 19558
rect 13436 19556 13460 19558
rect 13516 19556 13522 19558
rect 13214 19547 13522 19556
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9508 18034 9536 18090
rect 9324 16658 9352 18022
rect 9508 18006 9812 18034
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9600 16658 9628 16934
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 16250 8984 16390
rect 9692 16250 9720 16458
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 8852 16176 8904 16182
rect 8852 16118 8904 16124
rect 8864 15434 8892 16118
rect 9784 16114 9812 18006
rect 10214 17980 10522 17989
rect 10214 17978 10220 17980
rect 10276 17978 10300 17980
rect 10356 17978 10380 17980
rect 10436 17978 10460 17980
rect 10516 17978 10522 17980
rect 10276 17926 10278 17978
rect 10458 17926 10460 17978
rect 10214 17924 10220 17926
rect 10276 17924 10300 17926
rect 10356 17924 10380 17926
rect 10436 17924 10460 17926
rect 10516 17924 10522 17926
rect 10214 17915 10522 17924
rect 11532 17678 11560 18770
rect 12360 18766 12388 19382
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13004 18358 13032 18566
rect 12992 18352 13044 18358
rect 12992 18294 13044 18300
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 12544 17610 12572 18022
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11440 17270 11468 17478
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10152 16794 10180 17070
rect 10214 16892 10522 16901
rect 10214 16890 10220 16892
rect 10276 16890 10300 16892
rect 10356 16890 10380 16892
rect 10436 16890 10460 16892
rect 10516 16890 10522 16892
rect 10276 16838 10278 16890
rect 10458 16838 10460 16890
rect 10214 16836 10220 16838
rect 10276 16836 10300 16838
rect 10356 16836 10380 16838
rect 10436 16836 10460 16838
rect 10516 16836 10522 16838
rect 10214 16827 10522 16836
rect 10888 16794 10916 17070
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10152 16250 10180 16730
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 9784 15162 9812 16050
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 8956 14482 8984 14758
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13938 8800 14214
rect 9324 14074 9352 14282
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9692 14006 9720 14758
rect 9876 14346 9904 15370
rect 10152 14890 10180 16050
rect 10214 15804 10522 15813
rect 10214 15802 10220 15804
rect 10276 15802 10300 15804
rect 10356 15802 10380 15804
rect 10436 15802 10460 15804
rect 10516 15802 10522 15804
rect 10276 15750 10278 15802
rect 10458 15750 10460 15802
rect 10214 15748 10220 15750
rect 10276 15748 10300 15750
rect 10356 15748 10380 15750
rect 10436 15748 10460 15750
rect 10516 15748 10522 15750
rect 10214 15739 10522 15748
rect 10612 15026 10640 16730
rect 11440 16590 11468 17206
rect 11624 17202 11652 17478
rect 12544 17202 12572 17546
rect 12636 17202 12664 17818
rect 12900 17604 12952 17610
rect 12900 17546 12952 17552
rect 12912 17338 12940 17546
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 17338 13032 17478
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13096 17270 13124 19450
rect 13556 19174 13584 19774
rect 13648 19446 13676 19790
rect 14200 19514 14228 19790
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13214 18524 13522 18533
rect 13214 18522 13220 18524
rect 13276 18522 13300 18524
rect 13356 18522 13380 18524
rect 13436 18522 13460 18524
rect 13516 18522 13522 18524
rect 13276 18470 13278 18522
rect 13458 18470 13460 18522
rect 13214 18468 13220 18470
rect 13276 18468 13300 18470
rect 13356 18468 13380 18470
rect 13436 18468 13460 18470
rect 13516 18468 13522 18470
rect 13214 18459 13522 18468
rect 14292 18358 14320 20742
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13188 17610 13216 18022
rect 13464 17882 13492 18294
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13832 18170 13860 18226
rect 13740 18142 13860 18170
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13464 17610 13492 17818
rect 13740 17678 13768 18142
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 14292 17610 14320 18294
rect 13176 17604 13228 17610
rect 13176 17546 13228 17552
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 14280 17604 14332 17610
rect 14280 17546 14332 17552
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13214 17436 13522 17445
rect 13214 17434 13220 17436
rect 13276 17434 13300 17436
rect 13356 17434 13380 17436
rect 13436 17434 13460 17436
rect 13516 17434 13522 17436
rect 13276 17382 13278 17434
rect 13458 17382 13460 17434
rect 13214 17380 13220 17382
rect 13276 17380 13300 17382
rect 13356 17380 13380 17382
rect 13436 17380 13460 17382
rect 13516 17380 13522 17382
rect 13214 17371 13522 17380
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 13556 16998 13584 17478
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11164 15570 11192 16526
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11164 15026 11192 15506
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9692 13394 9720 13942
rect 9876 13410 9904 14282
rect 10060 13802 10088 14758
rect 10214 14716 10522 14725
rect 10214 14714 10220 14716
rect 10276 14714 10300 14716
rect 10356 14714 10380 14716
rect 10436 14714 10460 14716
rect 10516 14714 10522 14716
rect 10276 14662 10278 14714
rect 10458 14662 10460 14714
rect 10214 14660 10220 14662
rect 10276 14660 10300 14662
rect 10356 14660 10380 14662
rect 10436 14660 10460 14662
rect 10516 14660 10522 14662
rect 10214 14651 10522 14660
rect 10796 14618 10824 14962
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10612 13734 10640 14350
rect 11716 14074 11744 14962
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10214 13628 10522 13637
rect 10214 13626 10220 13628
rect 10276 13626 10300 13628
rect 10356 13626 10380 13628
rect 10436 13626 10460 13628
rect 10516 13626 10522 13628
rect 10276 13574 10278 13626
rect 10458 13574 10460 13626
rect 10214 13572 10220 13574
rect 10276 13572 10300 13574
rect 10356 13572 10380 13574
rect 10436 13572 10460 13574
rect 10516 13572 10522 13574
rect 10214 13563 10522 13572
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9784 13382 9904 13410
rect 10612 13394 10640 13670
rect 9956 13388 10008 13394
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8956 12434 8984 13126
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 8392 12378 8444 12384
rect 8496 12406 8616 12434
rect 8772 12406 8984 12434
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 10606 8432 11494
rect 8496 11082 8524 12406
rect 8772 12238 8800 12406
rect 9140 12238 9168 12922
rect 9324 12442 9352 13194
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8680 10266 8708 11698
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8956 11218 8984 11630
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9048 10810 9076 11222
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 9140 9994 9168 12174
rect 9416 11082 9444 12786
rect 9508 12782 9536 13262
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10742 9444 11018
rect 9404 10736 9456 10742
rect 9404 10678 9456 10684
rect 9508 10282 9536 12718
rect 9692 12434 9720 13330
rect 9784 13258 9812 13382
rect 9956 13330 10008 13336
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9784 12782 9812 13194
rect 9876 12986 9904 13262
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9968 12918 9996 13330
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12986 10916 13194
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 11900 12850 11928 16458
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15706 12480 15846
rect 12544 15706 12572 16390
rect 13214 16348 13522 16357
rect 13214 16346 13220 16348
rect 13276 16346 13300 16348
rect 13356 16346 13380 16348
rect 13436 16346 13460 16348
rect 13516 16346 13522 16348
rect 13276 16294 13278 16346
rect 13458 16294 13460 16346
rect 13214 16292 13220 16294
rect 13276 16292 13300 16294
rect 13356 16292 13380 16294
rect 13436 16292 13460 16294
rect 13516 16292 13522 16294
rect 13214 16283 13522 16292
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 15094 12572 15302
rect 12728 15162 12756 15438
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 14618 12480 14962
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12544 14414 12572 15030
rect 12820 14482 12848 15982
rect 13004 15638 13032 16050
rect 13648 15706 13676 17206
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16794 13768 16934
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13924 15706 13952 17138
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16590 14136 16934
rect 14292 16658 14320 17546
rect 14476 17202 14504 19654
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14108 15706 14136 15846
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 12992 15632 13044 15638
rect 12992 15574 13044 15580
rect 13004 15162 13032 15574
rect 14384 15502 14412 15846
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13096 15094 13124 15438
rect 13214 15260 13522 15269
rect 13214 15258 13220 15260
rect 13276 15258 13300 15260
rect 13356 15258 13380 15260
rect 13436 15258 13460 15260
rect 13516 15258 13522 15260
rect 13276 15206 13278 15258
rect 13458 15206 13460 15258
rect 13214 15204 13220 15206
rect 13276 15204 13300 15206
rect 13356 15204 13380 15206
rect 13436 15204 13460 15206
rect 13516 15204 13522 15206
rect 13214 15195 13522 15204
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 14200 14958 14228 15438
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14200 14482 14228 14894
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12820 14074 12848 14418
rect 13214 14172 13522 14181
rect 13214 14170 13220 14172
rect 13276 14170 13300 14172
rect 13356 14170 13380 14172
rect 13436 14170 13460 14172
rect 13516 14170 13522 14172
rect 13276 14118 13278 14170
rect 13458 14118 13460 14170
rect 13214 14116 13220 14118
rect 13276 14116 13300 14118
rect 13356 14116 13380 14118
rect 13436 14116 13460 14118
rect 13516 14116 13522 14118
rect 13214 14107 13522 14116
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 14200 13394 14228 14418
rect 14568 14006 14596 20810
rect 16132 20398 16160 20878
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 14740 20256 14792 20262
rect 15384 20256 15436 20262
rect 14740 20198 14792 20204
rect 15304 20216 15384 20244
rect 14752 20058 14780 20198
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 15304 19854 15332 20216
rect 15384 20198 15436 20204
rect 16214 20156 16522 20165
rect 16214 20154 16220 20156
rect 16276 20154 16300 20156
rect 16356 20154 16380 20156
rect 16436 20154 16460 20156
rect 16516 20154 16522 20156
rect 16276 20102 16278 20154
rect 16458 20102 16460 20154
rect 16214 20100 16220 20102
rect 16276 20100 16300 20102
rect 16356 20100 16380 20102
rect 16436 20100 16460 20102
rect 16516 20100 16522 20102
rect 16214 20091 16522 20100
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15304 18766 15332 19790
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16214 19068 16522 19077
rect 16214 19066 16220 19068
rect 16276 19066 16300 19068
rect 16356 19066 16380 19068
rect 16436 19066 16460 19068
rect 16516 19066 16522 19068
rect 16276 19014 16278 19066
rect 16458 19014 16460 19066
rect 16214 19012 16220 19014
rect 16276 19012 16300 19014
rect 16356 19012 16380 19014
rect 16436 19012 16460 19014
rect 16516 19012 16522 19014
rect 16214 19003 16522 19012
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15488 18086 15516 18634
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 17882 15516 18022
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15856 17678 15884 18294
rect 16132 17746 16160 18566
rect 16214 17980 16522 17989
rect 16214 17978 16220 17980
rect 16276 17978 16300 17980
rect 16356 17978 16380 17980
rect 16436 17978 16460 17980
rect 16516 17978 16522 17980
rect 16276 17926 16278 17978
rect 16458 17926 16460 17978
rect 16214 17924 16220 17926
rect 16276 17924 16300 17926
rect 16356 17924 16380 17926
rect 16436 17924 16460 17926
rect 16516 17924 16522 17926
rect 16214 17915 16522 17924
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 16214 16892 16522 16901
rect 16214 16890 16220 16892
rect 16276 16890 16300 16892
rect 16356 16890 16380 16892
rect 16436 16890 16460 16892
rect 16516 16890 16522 16892
rect 16276 16838 16278 16890
rect 16458 16838 16460 16890
rect 16214 16836 16220 16838
rect 16276 16836 16300 16838
rect 16356 16836 16380 16838
rect 16436 16836 16460 16838
rect 16516 16836 16522 16838
rect 16214 16827 16522 16836
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 14924 16448 14976 16454
rect 14976 16396 15056 16402
rect 14924 16390 15056 16396
rect 14936 16374 15056 16390
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 15028 15994 15056 16374
rect 15120 16250 15148 16594
rect 15488 16250 15516 16594
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 14660 15434 14688 15982
rect 15028 15966 15424 15994
rect 15396 15910 15424 15966
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 14648 15428 14700 15434
rect 14648 15370 14700 15376
rect 14660 15094 14688 15370
rect 14648 15088 14700 15094
rect 14648 15030 14700 15036
rect 15304 14482 15332 15846
rect 15580 15706 15608 16594
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15568 15700 15620 15706
rect 15568 15642 15620 15648
rect 15672 15366 15700 16050
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16132 15706 16160 15914
rect 16214 15804 16522 15813
rect 16214 15802 16220 15804
rect 16276 15802 16300 15804
rect 16356 15802 16380 15804
rect 16436 15802 16460 15804
rect 16516 15802 16522 15804
rect 16276 15750 16278 15802
rect 16458 15750 16460 15802
rect 16214 15748 16220 15750
rect 16276 15748 16300 15750
rect 16356 15748 16380 15750
rect 16436 15748 16460 15750
rect 16516 15748 16522 15750
rect 16214 15739 16522 15748
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15672 15162 15700 15302
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 16214 14716 16522 14725
rect 16214 14714 16220 14716
rect 16276 14714 16300 14716
rect 16356 14714 16380 14716
rect 16436 14714 16460 14716
rect 16516 14714 16522 14716
rect 16276 14662 16278 14714
rect 16458 14662 16460 14714
rect 16214 14660 16220 14662
rect 16276 14660 16300 14662
rect 16356 14660 16380 14662
rect 16436 14660 16460 14662
rect 16516 14660 16522 14662
rect 16214 14651 16522 14660
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 15672 13462 15700 14282
rect 16592 14074 16620 19382
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16684 18426 16712 19246
rect 16776 18970 16804 20402
rect 17052 19786 17080 20742
rect 17144 20262 17172 20810
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17880 20602 17908 20742
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17132 20256 17184 20262
rect 17132 20198 17184 20204
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16868 18970 16896 19110
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16776 18290 16804 18906
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16960 17678 16988 19450
rect 17052 18766 17080 19722
rect 17144 19718 17172 20198
rect 17328 19854 17356 20402
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17972 19854 18000 20198
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17132 19712 17184 19718
rect 17328 19666 17356 19790
rect 17132 19654 17184 19660
rect 17144 18970 17172 19654
rect 17236 19638 17356 19666
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17236 18766 17264 19638
rect 17420 18766 17448 19654
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17512 18086 17540 19654
rect 17696 18766 17724 19654
rect 17972 19174 18000 19790
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17972 18698 18000 19110
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17972 18154 18000 18634
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17500 18080 17552 18086
rect 17500 18022 17552 18028
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17604 16658 17632 18022
rect 18064 17882 18092 19314
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17038 15736 17094 15745
rect 17038 15671 17094 15680
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16684 14278 16712 14418
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15660 13456 15712 13462
rect 15660 13398 15712 13404
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12084 12986 12112 13126
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 9600 12406 9720 12434
rect 9600 12238 9628 12406
rect 10152 12238 10180 12582
rect 10214 12540 10522 12549
rect 10214 12538 10220 12540
rect 10276 12538 10300 12540
rect 10356 12538 10380 12540
rect 10436 12538 10460 12540
rect 10516 12538 10522 12540
rect 10276 12486 10278 12538
rect 10458 12486 10460 12538
rect 10214 12484 10220 12486
rect 10276 12484 10300 12486
rect 10356 12484 10380 12486
rect 10436 12484 10460 12486
rect 10516 12484 10522 12486
rect 10214 12475 10522 12484
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 11354 9812 11698
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9876 10538 9904 11494
rect 10214 11452 10522 11461
rect 10214 11450 10220 11452
rect 10276 11450 10300 11452
rect 10356 11450 10380 11452
rect 10436 11450 10460 11452
rect 10516 11450 10522 11452
rect 10276 11398 10278 11450
rect 10458 11398 10460 11450
rect 10214 11396 10220 11398
rect 10276 11396 10300 11398
rect 10356 11396 10380 11398
rect 10436 11396 10460 11398
rect 10516 11396 10522 11398
rect 10214 11387 10522 11396
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9508 10254 9628 10282
rect 9692 10266 9720 10406
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 7478 8432 8230
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8404 7002 8432 7414
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8496 6798 8524 7754
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8404 6458 8432 6666
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8024 5636 8076 5642
rect 8024 5578 8076 5584
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 7214 5468 7522 5477
rect 7214 5466 7220 5468
rect 7276 5466 7300 5468
rect 7356 5466 7380 5468
rect 7436 5466 7460 5468
rect 7516 5466 7522 5468
rect 7276 5414 7278 5466
rect 7458 5414 7460 5466
rect 7214 5412 7220 5414
rect 7276 5412 7300 5414
rect 7356 5412 7380 5414
rect 7436 5412 7460 5414
rect 7516 5412 7522 5414
rect 7214 5403 7522 5412
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6472 4826 6500 5102
rect 8220 5030 8248 5170
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 4160 4616 4212 4622
rect 4080 4576 4160 4604
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3804 4010 3832 4490
rect 4080 4434 4108 4576
rect 4160 4558 4212 4564
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 3988 4406 4108 4434
rect 3792 4004 3844 4010
rect 3792 3946 3844 3952
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3804 2854 3832 3946
rect 3988 3738 4016 4406
rect 7214 4380 7522 4389
rect 7214 4378 7220 4380
rect 7276 4378 7300 4380
rect 7356 4378 7380 4380
rect 7436 4378 7460 4380
rect 7516 4378 7522 4380
rect 7276 4326 7278 4378
rect 7458 4326 7460 4378
rect 7214 4324 7220 4326
rect 7276 4324 7300 4326
rect 7356 4324 7380 4326
rect 7436 4324 7460 4326
rect 7516 4324 7522 4326
rect 7214 4315 7522 4324
rect 8220 4128 8248 4966
rect 8312 4622 8340 5238
rect 8404 4622 8432 5510
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4146 8432 4422
rect 8496 4146 8524 4490
rect 8300 4140 8352 4146
rect 8220 4100 8300 4128
rect 8300 4082 8352 4088
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 4080 3738 4108 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 7024 3534 7052 3878
rect 8036 3602 8064 3878
rect 8312 3602 8340 4082
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 4356 3126 4384 3470
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5460 3194 5488 3402
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7024 2514 7052 3470
rect 7214 3292 7522 3301
rect 7214 3290 7220 3292
rect 7276 3290 7300 3292
rect 7356 3290 7380 3292
rect 7436 3290 7460 3292
rect 7516 3290 7522 3292
rect 7276 3238 7278 3290
rect 7458 3238 7460 3290
rect 7214 3236 7220 3238
rect 7276 3236 7300 3238
rect 7356 3236 7380 3238
rect 7436 3236 7460 3238
rect 7516 3236 7522 3238
rect 7214 3227 7522 3236
rect 8404 3194 8432 4082
rect 8588 3534 8616 9318
rect 8772 8906 8800 9930
rect 9600 9704 9628 10254
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9784 9722 9812 10202
rect 9968 9994 9996 10406
rect 10060 10266 10088 10406
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9048 9676 9628 9704
rect 9048 9586 9076 9676
rect 9600 9586 9628 9676
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8772 8566 8800 8842
rect 9048 8838 9076 9386
rect 9140 9178 9168 9522
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 9178 9260 9318
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9324 8634 9352 9386
rect 9876 9024 9904 9658
rect 9692 8996 9904 9024
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9416 8566 9444 8910
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8864 7954 8892 8434
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8864 6798 8892 7890
rect 9416 7546 9444 8502
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9692 6338 9720 8996
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9784 6866 9812 8842
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9876 7002 9904 8230
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9416 6310 9720 6338
rect 9772 6316 9824 6322
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5370 8708 6054
rect 9416 5914 9444 6310
rect 9772 6258 9824 6264
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8772 5234 8800 5646
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8852 5228 8904 5234
rect 8852 5170 8904 5176
rect 8772 4486 8800 5170
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8864 4146 8892 5170
rect 9140 4758 9168 5646
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9324 5302 9352 5510
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9416 5234 9444 5510
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9140 4282 9168 4694
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9232 4162 9260 4490
rect 9232 4146 9352 4162
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9220 4140 9352 4146
rect 9272 4134 9352 4140
rect 9220 4082 9272 4088
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8864 3738 8892 3878
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 9140 3534 9168 4082
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9232 3534 9260 3946
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8956 3058 8984 3334
rect 9232 3194 9260 3470
rect 9324 3466 9352 4134
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9416 3126 9444 5170
rect 9508 4010 9536 6190
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5370 9720 5578
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9784 4486 9812 6258
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9600 3534 9628 4082
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3738 9720 3878
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 9784 2446 9812 4422
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9968 3194 9996 3334
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10060 2582 10088 9862
rect 10152 9586 10180 10610
rect 10214 10364 10522 10373
rect 10214 10362 10220 10364
rect 10276 10362 10300 10364
rect 10356 10362 10380 10364
rect 10436 10362 10460 10364
rect 10516 10362 10522 10364
rect 10276 10310 10278 10362
rect 10458 10310 10460 10362
rect 10214 10308 10220 10310
rect 10276 10308 10300 10310
rect 10356 10308 10380 10310
rect 10436 10308 10460 10310
rect 10516 10308 10522 10310
rect 10214 10299 10522 10308
rect 10612 10266 10640 11154
rect 10888 11150 10916 11494
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10704 10062 10732 10610
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10152 9042 10180 9522
rect 10214 9276 10522 9285
rect 10214 9274 10220 9276
rect 10276 9274 10300 9276
rect 10356 9274 10380 9276
rect 10436 9274 10460 9276
rect 10516 9274 10522 9276
rect 10276 9222 10278 9274
rect 10458 9222 10460 9274
rect 10214 9220 10220 9222
rect 10276 9220 10300 9222
rect 10356 9220 10380 9222
rect 10436 9220 10460 9222
rect 10516 9220 10522 9222
rect 10214 9211 10522 9220
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10152 8362 10180 8978
rect 10520 8566 10548 8978
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10214 8188 10522 8197
rect 10214 8186 10220 8188
rect 10276 8186 10300 8188
rect 10356 8186 10380 8188
rect 10436 8186 10460 8188
rect 10516 8186 10522 8188
rect 10276 8134 10278 8186
rect 10458 8134 10460 8186
rect 10214 8132 10220 8134
rect 10276 8132 10300 8134
rect 10356 8132 10380 8134
rect 10436 8132 10460 8134
rect 10516 8132 10522 8134
rect 10214 8123 10522 8132
rect 10612 8090 10640 9998
rect 10796 9722 10824 10406
rect 10888 10130 10916 10610
rect 11072 10470 11100 11018
rect 11164 10674 11192 11630
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 11072 9042 11100 10406
rect 11348 10062 11376 10678
rect 12176 10606 12204 13194
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13096 12850 13124 13126
rect 13214 13084 13522 13093
rect 13214 13082 13220 13084
rect 13276 13082 13300 13084
rect 13356 13082 13380 13084
rect 13436 13082 13460 13084
rect 13516 13082 13522 13084
rect 13276 13030 13278 13082
rect 13458 13030 13460 13082
rect 13214 13028 13220 13030
rect 13276 13028 13300 13030
rect 13356 13028 13380 13030
rect 13436 13028 13460 13030
rect 13516 13028 13522 13030
rect 13214 13019 13522 13028
rect 13648 12986 13676 13126
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 12452 9722 12480 10610
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12544 9586 12572 12038
rect 12728 11354 12756 12174
rect 13096 11898 13124 12786
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13214 11996 13522 12005
rect 13214 11994 13220 11996
rect 13276 11994 13300 11996
rect 13356 11994 13380 11996
rect 13436 11994 13460 11996
rect 13516 11994 13522 11996
rect 13276 11942 13278 11994
rect 13458 11942 13460 11994
rect 13214 11940 13220 11942
rect 13276 11940 13300 11942
rect 13356 11940 13380 11942
rect 13436 11940 13460 11942
rect 13516 11940 13522 11942
rect 13214 11931 13522 11940
rect 13648 11898 13676 12718
rect 13740 12646 13768 13126
rect 14568 12986 14596 13194
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12442 13768 12582
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 14108 12238 14136 12922
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15304 12646 15332 12854
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15580 12238 15608 12718
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 14384 11830 14412 12174
rect 15672 12102 15700 12650
rect 15764 12434 15792 13874
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16214 13628 16522 13637
rect 16214 13626 16220 13628
rect 16276 13626 16300 13628
rect 16356 13626 16380 13628
rect 16436 13626 16460 13628
rect 16516 13626 16522 13628
rect 16276 13574 16278 13626
rect 16458 13574 16460 13626
rect 16214 13572 16220 13574
rect 16276 13572 16300 13574
rect 16356 13572 16380 13574
rect 16436 13572 16460 13574
rect 16516 13572 16522 13574
rect 16214 13563 16522 13572
rect 16592 13462 16620 13670
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16040 12986 16068 13126
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16316 12918 16344 13126
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16214 12540 16522 12549
rect 16214 12538 16220 12540
rect 16276 12538 16300 12540
rect 16356 12538 16380 12540
rect 16436 12538 16460 12540
rect 16516 12538 16522 12540
rect 16276 12486 16278 12538
rect 16458 12486 16460 12538
rect 16214 12484 16220 12486
rect 16276 12484 16300 12486
rect 16356 12484 16380 12486
rect 16436 12484 16460 12486
rect 16516 12484 16522 12486
rect 16214 12475 16522 12484
rect 16592 12434 16620 13262
rect 16684 13190 16712 14214
rect 17052 13530 17080 15671
rect 17328 15502 17356 16594
rect 17696 16590 17724 17478
rect 17972 17270 18000 17682
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17972 16590 18000 17206
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 18064 16522 18092 17546
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 17604 15502 17632 16458
rect 18156 16114 18184 16934
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 15502 17908 15846
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 13734 17172 14350
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 17144 12986 17172 13670
rect 16672 12980 16724 12986
rect 17132 12980 17184 12986
rect 16724 12940 16896 12968
rect 16672 12922 16724 12928
rect 15764 12406 15884 12434
rect 16592 12406 16804 12434
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 14372 11824 14424 11830
rect 15856 11778 15884 12406
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15948 11830 15976 12106
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 14372 11766 14424 11772
rect 14384 11558 14412 11766
rect 15764 11762 15884 11778
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 15752 11756 15884 11762
rect 15804 11750 15884 11756
rect 15752 11698 15804 11704
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12636 10742 12664 10950
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 13096 10470 13124 10950
rect 13214 10908 13522 10917
rect 13214 10906 13220 10908
rect 13276 10906 13300 10908
rect 13356 10906 13380 10908
rect 13436 10906 13460 10908
rect 13516 10906 13522 10908
rect 13276 10854 13278 10906
rect 13458 10854 13460 10906
rect 13214 10852 13220 10854
rect 13276 10852 13300 10854
rect 13356 10852 13380 10854
rect 13436 10852 13460 10854
rect 13516 10852 13522 10854
rect 13214 10843 13522 10852
rect 13832 10674 13860 11018
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10784 8900 10836 8906
rect 10784 8842 10836 8848
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10704 8022 10732 8434
rect 10796 8090 10824 8842
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10692 8016 10744 8022
rect 10692 7958 10744 7964
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10704 7410 10732 7686
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10508 7268 10560 7274
rect 10796 7256 10824 7754
rect 10888 7410 10916 7958
rect 10980 7562 11008 8434
rect 11164 7698 11192 8774
rect 11256 8022 11284 9318
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11244 8016 11296 8022
rect 11244 7958 11296 7964
rect 11164 7670 11284 7698
rect 10980 7534 11192 7562
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10560 7228 10824 7256
rect 10508 7210 10560 7216
rect 10214 7100 10522 7109
rect 10214 7098 10220 7100
rect 10276 7098 10300 7100
rect 10356 7098 10380 7100
rect 10436 7098 10460 7100
rect 10516 7098 10522 7100
rect 10276 7046 10278 7098
rect 10458 7046 10460 7098
rect 10214 7044 10220 7046
rect 10276 7044 10300 7046
rect 10356 7044 10380 7046
rect 10436 7044 10460 7046
rect 10516 7044 10522 7046
rect 10214 7035 10522 7044
rect 10796 6730 10824 7228
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10888 6798 10916 7210
rect 10980 7002 11008 7346
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11164 6798 11192 7534
rect 11256 7342 11284 7670
rect 11348 7478 11376 8842
rect 11624 8430 11652 9318
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11428 8424 11480 8430
rect 11612 8424 11664 8430
rect 11428 8366 11480 8372
rect 11532 8384 11612 8412
rect 11440 7886 11468 8366
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11428 7744 11480 7750
rect 11532 7732 11560 8384
rect 11612 8366 11664 8372
rect 11480 7704 11560 7732
rect 11428 7686 11480 7692
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6338 10824 6666
rect 10796 6310 10916 6338
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 10152 5914 10180 6122
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10214 6012 10522 6021
rect 10214 6010 10220 6012
rect 10276 6010 10300 6012
rect 10356 6010 10380 6012
rect 10436 6010 10460 6012
rect 10516 6010 10522 6012
rect 10276 5958 10278 6010
rect 10458 5958 10460 6010
rect 10214 5956 10220 5958
rect 10276 5956 10300 5958
rect 10356 5956 10380 5958
rect 10436 5956 10460 5958
rect 10516 5956 10522 5958
rect 10214 5947 10522 5956
rect 10796 5914 10824 6054
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10888 5710 10916 6310
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10214 4924 10522 4933
rect 10214 4922 10220 4924
rect 10276 4922 10300 4924
rect 10356 4922 10380 4924
rect 10436 4922 10460 4924
rect 10516 4922 10522 4924
rect 10276 4870 10278 4922
rect 10458 4870 10460 4922
rect 10214 4868 10220 4870
rect 10276 4868 10300 4870
rect 10356 4868 10380 4870
rect 10436 4868 10460 4870
rect 10516 4868 10522 4870
rect 10214 4859 10522 4868
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10214 3836 10522 3845
rect 10214 3834 10220 3836
rect 10276 3834 10300 3836
rect 10356 3834 10380 3836
rect 10436 3834 10460 3836
rect 10516 3834 10522 3836
rect 10276 3782 10278 3834
rect 10458 3782 10460 3834
rect 10214 3780 10220 3782
rect 10276 3780 10300 3782
rect 10356 3780 10380 3782
rect 10436 3780 10460 3782
rect 10516 3780 10522 3782
rect 10214 3771 10522 3780
rect 10416 2984 10468 2990
rect 10468 2944 10640 2972
rect 10416 2926 10468 2932
rect 10214 2748 10522 2757
rect 10214 2746 10220 2748
rect 10276 2746 10300 2748
rect 10356 2746 10380 2748
rect 10436 2746 10460 2748
rect 10516 2746 10522 2748
rect 10276 2694 10278 2746
rect 10458 2694 10460 2746
rect 10214 2692 10220 2694
rect 10276 2692 10300 2694
rect 10356 2692 10380 2694
rect 10436 2692 10460 2694
rect 10516 2692 10522 2694
rect 10214 2683 10522 2692
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 5276 1306 5304 2382
rect 7214 2204 7522 2213
rect 7214 2202 7220 2204
rect 7276 2202 7300 2204
rect 7356 2202 7380 2204
rect 7436 2202 7460 2204
rect 7516 2202 7522 2204
rect 7276 2150 7278 2202
rect 7458 2150 7460 2202
rect 7214 2148 7220 2150
rect 7276 2148 7300 2150
rect 7356 2148 7380 2150
rect 7436 2148 7460 2150
rect 7516 2148 7522 2150
rect 7214 2139 7522 2148
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 10336 870 10456 898
rect 10336 800 10364 870
rect 18 0 74 800
rect 5170 0 5226 800
rect 10322 0 10378 800
rect 10428 762 10456 870
rect 10612 762 10640 2944
rect 10888 2446 10916 4490
rect 10980 4146 11008 6258
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11164 5302 11192 5510
rect 11348 5302 11376 7414
rect 11808 7274 11836 8910
rect 12164 8900 12216 8906
rect 12164 8842 12216 8848
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11900 7546 11928 7822
rect 12084 7818 12112 8774
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11796 7268 11848 7274
rect 11796 7210 11848 7216
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5574 11560 6054
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4214 11100 4966
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 2650 11008 4082
rect 11256 2650 11284 5170
rect 11716 4826 11744 6258
rect 12176 6254 12204 8842
rect 12452 8566 12480 8978
rect 12636 8634 12664 9522
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 8634 12848 8774
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 7954 12296 8230
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12360 5914 12388 6258
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 12452 3738 12480 8502
rect 13096 8294 13124 10406
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13214 9820 13522 9829
rect 13214 9818 13220 9820
rect 13276 9818 13300 9820
rect 13356 9818 13380 9820
rect 13436 9818 13460 9820
rect 13516 9818 13522 9820
rect 13276 9766 13278 9818
rect 13458 9766 13460 9818
rect 13214 9764 13220 9766
rect 13276 9764 13300 9766
rect 13356 9764 13380 9766
rect 13436 9764 13460 9766
rect 13516 9764 13522 9766
rect 13214 9755 13522 9764
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13214 8732 13522 8741
rect 13214 8730 13220 8732
rect 13276 8730 13300 8732
rect 13356 8730 13380 8732
rect 13436 8730 13460 8732
rect 13516 8730 13522 8732
rect 13276 8678 13278 8730
rect 13458 8678 13460 8730
rect 13214 8676 13220 8678
rect 13276 8676 13300 8678
rect 13356 8676 13380 8678
rect 13436 8676 13460 8678
rect 13516 8676 13522 8678
rect 13214 8667 13522 8676
rect 13556 8634 13584 8774
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 13556 7818 13584 8434
rect 13832 8430 13860 9998
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 13214 7644 13522 7653
rect 13214 7642 13220 7644
rect 13276 7642 13300 7644
rect 13356 7642 13380 7644
rect 13436 7642 13460 7644
rect 13516 7642 13522 7644
rect 13276 7590 13278 7642
rect 13458 7590 13460 7642
rect 13214 7588 13220 7590
rect 13276 7588 13300 7590
rect 13356 7588 13380 7590
rect 13436 7588 13460 7590
rect 13516 7588 13522 7590
rect 13214 7579 13522 7588
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12544 5166 12572 6190
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12544 4282 12572 5102
rect 12636 4622 12664 5510
rect 12820 5370 12848 7346
rect 13214 6556 13522 6565
rect 13214 6554 13220 6556
rect 13276 6554 13300 6556
rect 13356 6554 13380 6556
rect 13436 6554 13460 6556
rect 13516 6554 13522 6556
rect 13276 6502 13278 6554
rect 13458 6502 13460 6554
rect 13214 6500 13220 6502
rect 13276 6500 13300 6502
rect 13356 6500 13380 6502
rect 13436 6500 13460 6502
rect 13516 6500 13522 6502
rect 13214 6491 13522 6500
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13556 5710 13584 5782
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13214 5468 13522 5477
rect 13214 5466 13220 5468
rect 13276 5466 13300 5468
rect 13356 5466 13380 5468
rect 13436 5466 13460 5468
rect 13516 5466 13522 5468
rect 13276 5414 13278 5466
rect 13458 5414 13460 5466
rect 13214 5412 13220 5414
rect 13276 5412 13300 5414
rect 13356 5412 13380 5414
rect 13436 5412 13460 5414
rect 13516 5412 13522 5414
rect 13214 5403 13522 5412
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13280 4826 13308 5034
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13372 4826 13400 4966
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 13556 4486 13584 5646
rect 13924 5302 13952 11154
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14200 10266 14228 10542
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14384 10062 14412 11494
rect 15856 11082 15884 11750
rect 15948 11150 15976 11766
rect 16684 11558 16712 12038
rect 16776 11898 16804 12406
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16764 11620 16816 11626
rect 16764 11562 16816 11568
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16214 11452 16522 11461
rect 16214 11450 16220 11452
rect 16276 11450 16300 11452
rect 16356 11450 16380 11452
rect 16436 11450 16460 11452
rect 16516 11450 16522 11452
rect 16276 11398 16278 11450
rect 16458 11398 16460 11450
rect 16214 11396 16220 11398
rect 16276 11396 16300 11398
rect 16356 11396 16380 11398
rect 16436 11396 16460 11398
rect 16516 11396 16522 11398
rect 16214 11387 16522 11396
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14384 9586 14412 9998
rect 14648 9988 14700 9994
rect 14648 9930 14700 9936
rect 14660 9654 14688 9930
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 15212 9382 15240 10678
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14292 7818 14320 8570
rect 15396 8294 15424 8774
rect 15856 8498 15884 11018
rect 15948 10266 15976 11086
rect 16776 11082 16804 11562
rect 16868 11558 16896 12940
rect 17132 12922 17184 12928
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 17144 11558 17172 12650
rect 17328 11762 17356 14214
rect 17420 13530 17448 14554
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 12968 17724 13262
rect 17604 12940 17724 12968
rect 17604 12306 17632 12940
rect 17880 12918 17908 13466
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17236 11354 17264 11630
rect 17604 11354 17632 12242
rect 17972 11830 18000 15370
rect 18156 15026 18184 16050
rect 18248 15638 18276 21286
rect 19214 20700 19522 20709
rect 19214 20698 19220 20700
rect 19276 20698 19300 20700
rect 19356 20698 19380 20700
rect 19436 20698 19460 20700
rect 19516 20698 19522 20700
rect 19276 20646 19278 20698
rect 19458 20646 19460 20698
rect 19214 20644 19220 20646
rect 19276 20644 19300 20646
rect 19356 20644 19380 20646
rect 19436 20644 19460 20646
rect 19516 20644 19522 20646
rect 19214 20635 19522 20644
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19812 19786 19840 20198
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19214 19612 19522 19621
rect 19214 19610 19220 19612
rect 19276 19610 19300 19612
rect 19356 19610 19380 19612
rect 19436 19610 19460 19612
rect 19516 19610 19522 19612
rect 19276 19558 19278 19610
rect 19458 19558 19460 19610
rect 19214 19556 19220 19558
rect 19276 19556 19300 19558
rect 19356 19556 19380 19558
rect 19436 19556 19460 19558
rect 19516 19556 19522 19558
rect 19214 19547 19522 19556
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18800 18970 18828 19314
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19214 18524 19522 18533
rect 19214 18522 19220 18524
rect 19276 18522 19300 18524
rect 19356 18522 19380 18524
rect 19436 18522 19460 18524
rect 19516 18522 19522 18524
rect 19276 18470 19278 18522
rect 19458 18470 19460 18522
rect 19214 18468 19220 18470
rect 19276 18468 19300 18470
rect 19356 18468 19380 18470
rect 19436 18468 19460 18470
rect 19516 18468 19522 18470
rect 19214 18459 19522 18468
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18616 16794 18644 17750
rect 19444 17678 19472 18294
rect 19628 17882 19656 18702
rect 19812 18630 19840 19722
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19904 18902 19932 19110
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19720 18426 19748 18566
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19214 17436 19522 17445
rect 19214 17434 19220 17436
rect 19276 17434 19300 17436
rect 19356 17434 19380 17436
rect 19436 17434 19460 17436
rect 19516 17434 19522 17436
rect 19276 17382 19278 17434
rect 19458 17382 19460 17434
rect 19214 17380 19220 17382
rect 19276 17380 19300 17382
rect 19356 17380 19380 17382
rect 19436 17380 19460 17382
rect 19516 17380 19522 17382
rect 19214 17371 19522 17380
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 18708 16794 18736 17138
rect 19628 16794 19656 17138
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 18984 16182 19012 16458
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18236 15632 18288 15638
rect 18236 15574 18288 15580
rect 18236 15360 18288 15366
rect 18236 15302 18288 15308
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18156 14414 18184 14962
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18156 14074 18184 14350
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13326 18092 13806
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18064 12850 18092 13262
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 18064 11898 18092 12106
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 18156 11506 18184 12038
rect 17880 11478 18184 11506
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16776 10810 16804 11018
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16214 10364 16522 10373
rect 16214 10362 16220 10364
rect 16276 10362 16300 10364
rect 16356 10362 16380 10364
rect 16436 10362 16460 10364
rect 16516 10362 16522 10364
rect 16276 10310 16278 10362
rect 16458 10310 16460 10362
rect 16214 10308 16220 10310
rect 16276 10308 16300 10310
rect 16356 10308 16380 10310
rect 16436 10308 16460 10310
rect 16516 10308 16522 10310
rect 16214 10299 16522 10308
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5914 14228 6054
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12544 3618 12572 4218
rect 12912 4146 12940 4422
rect 13214 4380 13522 4389
rect 13214 4378 13220 4380
rect 13276 4378 13300 4380
rect 13356 4378 13380 4380
rect 13436 4378 13460 4380
rect 13516 4378 13522 4380
rect 13276 4326 13278 4378
rect 13458 4326 13460 4378
rect 13214 4324 13220 4326
rect 13276 4324 13300 4326
rect 13356 4324 13380 4326
rect 13436 4324 13460 4326
rect 13516 4324 13522 4326
rect 13214 4315 13522 4324
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12452 3590 12572 3618
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 11532 3194 11560 3402
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11808 2446 11836 3334
rect 12452 3058 12480 3590
rect 12820 3534 12848 3878
rect 13556 3670 13584 4422
rect 13740 4282 13768 4422
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13832 3738 13860 4558
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 12808 3528 12860 3534
rect 12728 3488 12808 3516
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12544 3058 12572 3402
rect 12728 3194 12756 3488
rect 12808 3470 12860 3476
rect 13214 3292 13522 3301
rect 13214 3290 13220 3292
rect 13276 3290 13300 3292
rect 13356 3290 13380 3292
rect 13436 3290 13460 3292
rect 13516 3290 13522 3292
rect 13276 3238 13278 3290
rect 13458 3238 13460 3290
rect 13214 3236 13220 3238
rect 13276 3236 13300 3238
rect 13356 3236 13380 3238
rect 13436 3236 13460 3238
rect 13516 3236 13522 3238
rect 13214 3227 13522 3236
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 2650 12112 2926
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12268 2446 12296 2994
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12360 2514 12388 2790
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12452 2446 12480 2994
rect 12544 2650 12572 2994
rect 13556 2854 13584 3606
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3194 13768 3334
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 14108 2582 14136 3470
rect 14292 3126 14320 7754
rect 15212 7018 15240 7822
rect 15396 7818 15424 8230
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15120 7002 15240 7018
rect 15120 6996 15252 7002
rect 15120 6990 15200 6996
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14384 5370 14412 6258
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14476 5370 14504 6190
rect 15120 5778 15148 6990
rect 15200 6938 15252 6944
rect 15488 6798 15516 7142
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15580 6730 15608 8298
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15856 5710 15884 8434
rect 15948 7478 15976 8502
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16040 8090 16068 8230
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 16132 7886 16160 9998
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16214 9276 16522 9285
rect 16214 9274 16220 9276
rect 16276 9274 16300 9276
rect 16356 9274 16380 9276
rect 16436 9274 16460 9276
rect 16516 9274 16522 9276
rect 16276 9222 16278 9274
rect 16458 9222 16460 9274
rect 16214 9220 16220 9222
rect 16276 9220 16300 9222
rect 16356 9220 16380 9222
rect 16436 9220 16460 9222
rect 16516 9220 16522 9222
rect 16214 9211 16522 9220
rect 16592 9042 16620 9318
rect 17788 9178 17816 11154
rect 17880 10674 17908 11478
rect 18156 11354 18184 11478
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18064 10674 18092 11290
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18248 10266 18276 15302
rect 19076 15094 19104 16458
rect 19628 16454 19656 16730
rect 19720 16590 19748 18022
rect 19812 17678 19840 18566
rect 19904 18358 19932 18838
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 19996 17746 20024 18634
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19214 16348 19522 16357
rect 19214 16346 19220 16348
rect 19276 16346 19300 16348
rect 19356 16346 19380 16348
rect 19436 16346 19460 16348
rect 19516 16346 19522 16348
rect 19276 16294 19278 16346
rect 19458 16294 19460 16346
rect 19214 16292 19220 16294
rect 19276 16292 19300 16294
rect 19356 16292 19380 16294
rect 19436 16292 19460 16294
rect 19516 16292 19522 16294
rect 19214 16283 19522 16292
rect 19628 16250 19656 16390
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19892 16176 19944 16182
rect 19892 16118 19944 16124
rect 19214 15260 19522 15269
rect 19214 15258 19220 15260
rect 19276 15258 19300 15260
rect 19356 15258 19380 15260
rect 19436 15258 19460 15260
rect 19516 15258 19522 15260
rect 19276 15206 19278 15258
rect 19458 15206 19460 15258
rect 19214 15204 19220 15206
rect 19276 15204 19300 15206
rect 19356 15204 19380 15206
rect 19436 15204 19460 15206
rect 19516 15204 19522 15206
rect 19214 15195 19522 15204
rect 19904 15162 19932 16118
rect 20272 15502 20300 21490
rect 20444 21344 20496 21350
rect 20444 21286 20496 21292
rect 20456 21185 20484 21286
rect 20442 21176 20498 21185
rect 20442 21111 20498 21120
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 18984 14006 19012 14214
rect 19214 14172 19522 14181
rect 19214 14170 19220 14172
rect 19276 14170 19300 14172
rect 19356 14170 19380 14172
rect 19436 14170 19460 14172
rect 19516 14170 19522 14172
rect 19276 14118 19278 14170
rect 19458 14118 19460 14170
rect 19214 14116 19220 14118
rect 19276 14116 19300 14118
rect 19356 14116 19380 14118
rect 19436 14116 19460 14118
rect 19516 14116 19522 14118
rect 19214 14107 19522 14116
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 18984 12918 19012 13942
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19214 13084 19522 13093
rect 19214 13082 19220 13084
rect 19276 13082 19300 13084
rect 19356 13082 19380 13084
rect 19436 13082 19460 13084
rect 19516 13082 19522 13084
rect 19276 13030 19278 13082
rect 19458 13030 19460 13082
rect 19214 13028 19220 13030
rect 19276 13028 19300 13030
rect 19356 13028 19380 13030
rect 19436 13028 19460 13030
rect 19516 13028 19522 13030
rect 19214 13019 19522 13028
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 18512 12912 18564 12918
rect 18512 12854 18564 12860
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18340 11762 18368 12582
rect 18524 12434 18552 12854
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18524 12406 18736 12434
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18616 11830 18644 12310
rect 18708 12238 18736 12406
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18800 12050 18828 12718
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 18892 12306 18920 12650
rect 19260 12442 19288 12922
rect 19996 12918 20024 13670
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 19260 12186 19288 12378
rect 19536 12374 19564 12786
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19076 12158 19288 12186
rect 20168 12164 20220 12170
rect 18800 12022 19012 12050
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18984 11762 19012 12022
rect 19076 11830 19104 12158
rect 20168 12106 20220 12112
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19214 11996 19522 12005
rect 19214 11994 19220 11996
rect 19276 11994 19300 11996
rect 19356 11994 19380 11996
rect 19436 11994 19460 11996
rect 19516 11994 19522 11996
rect 19276 11942 19278 11994
rect 19458 11942 19460 11994
rect 19214 11940 19220 11942
rect 19276 11940 19300 11942
rect 19356 11940 19380 11942
rect 19436 11940 19460 11942
rect 19516 11940 19522 11942
rect 19214 11931 19522 11940
rect 19904 11898 19932 12038
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 20180 11830 20208 12106
rect 19064 11824 19116 11830
rect 19064 11766 19116 11772
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19214 10908 19522 10917
rect 19214 10906 19220 10908
rect 19276 10906 19300 10908
rect 19356 10906 19380 10908
rect 19436 10906 19460 10908
rect 19516 10906 19522 10908
rect 19276 10854 19278 10906
rect 19458 10854 19460 10906
rect 19214 10852 19220 10854
rect 19276 10852 19300 10854
rect 19356 10852 19380 10854
rect 19436 10852 19460 10854
rect 19516 10852 19522 10854
rect 19214 10843 19522 10852
rect 19628 10810 19656 11290
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19616 10804 19668 10810
rect 19616 10746 19668 10752
rect 19720 10674 19748 11018
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18328 10056 18380 10062
rect 18064 10004 18328 10010
rect 18064 9998 18380 10004
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18064 9982 18368 9998
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 18064 9110 18092 9982
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18156 9178 18184 9862
rect 18248 9722 18276 9862
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 18144 9036 18196 9042
rect 18248 9024 18276 9658
rect 18708 9178 18736 9998
rect 18800 9722 18828 10610
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19628 10198 19656 10406
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19214 9820 19522 9829
rect 19214 9818 19220 9820
rect 19276 9818 19300 9820
rect 19356 9818 19380 9820
rect 19436 9818 19460 9820
rect 19516 9818 19522 9820
rect 19276 9766 19278 9818
rect 19458 9766 19460 9818
rect 19214 9764 19220 9766
rect 19276 9764 19300 9766
rect 19356 9764 19380 9766
rect 19436 9764 19460 9766
rect 19516 9764 19522 9766
rect 19214 9755 19522 9764
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 19720 9586 19748 10610
rect 19812 10538 19840 11086
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 20088 10674 20116 10950
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19800 10532 19852 10538
rect 19800 10474 19852 10480
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18196 8996 18276 9024
rect 18144 8978 18196 8984
rect 16592 8566 16620 8978
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16214 8188 16522 8197
rect 16214 8186 16220 8188
rect 16276 8186 16300 8188
rect 16356 8186 16380 8188
rect 16436 8186 16460 8188
rect 16516 8186 16522 8188
rect 16276 8134 16278 8186
rect 16458 8134 16460 8186
rect 16214 8132 16220 8134
rect 16276 8132 16300 8134
rect 16356 8132 16380 8134
rect 16436 8132 16460 8134
rect 16516 8132 16522 8134
rect 16214 8123 16522 8132
rect 16592 7886 16620 8502
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 16132 7410 16160 7822
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7478 16528 7686
rect 17236 7546 17264 8026
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16214 7100 16522 7109
rect 16214 7098 16220 7100
rect 16276 7098 16300 7100
rect 16356 7098 16380 7100
rect 16436 7098 16460 7100
rect 16516 7098 16522 7100
rect 16276 7046 16278 7098
rect 16458 7046 16460 7098
rect 16214 7044 16220 7046
rect 16276 7044 16300 7046
rect 16356 7044 16380 7046
rect 16436 7044 16460 7046
rect 16516 7044 16522 7046
rect 16214 7035 16522 7044
rect 16592 6662 16620 7278
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16960 6662 16988 7142
rect 17052 6934 17080 7346
rect 17040 6928 17092 6934
rect 17040 6870 17092 6876
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16214 6012 16522 6021
rect 16214 6010 16220 6012
rect 16276 6010 16300 6012
rect 16356 6010 16380 6012
rect 16436 6010 16460 6012
rect 16516 6010 16522 6012
rect 16276 5958 16278 6010
rect 16458 5958 16460 6010
rect 16214 5956 16220 5958
rect 16276 5956 16300 5958
rect 16356 5956 16380 5958
rect 16436 5956 16460 5958
rect 16516 5956 16522 5958
rect 16214 5947 16522 5956
rect 16592 5710 16620 6598
rect 16960 6322 16988 6598
rect 17052 6458 17080 6870
rect 17328 6866 17356 8774
rect 17604 8090 17632 8842
rect 17696 8498 17724 8910
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 18064 8634 18092 8842
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17696 7886 17724 8434
rect 18800 8090 18828 8774
rect 18984 8634 19012 9454
rect 19214 8732 19522 8741
rect 19214 8730 19220 8732
rect 19276 8730 19300 8732
rect 19356 8730 19380 8732
rect 19436 8730 19460 8732
rect 19516 8730 19522 8732
rect 19276 8678 19278 8730
rect 19458 8678 19460 8730
rect 19214 8676 19220 8678
rect 19276 8676 19300 8678
rect 19356 8676 19380 8678
rect 19436 8676 19460 8678
rect 19516 8676 19522 8678
rect 19214 8667 19522 8676
rect 19720 8634 19748 9522
rect 20088 9382 20116 10610
rect 20180 10266 20208 11766
rect 20810 10296 20866 10305
rect 20168 10260 20220 10266
rect 20810 10231 20866 10240
rect 20168 10202 20220 10208
rect 20180 10062 20208 10202
rect 20824 10062 20852 10231
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 19076 8022 19104 8434
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19064 8016 19116 8022
rect 19524 8016 19576 8022
rect 19116 7964 19524 7970
rect 19064 7958 19576 7964
rect 19076 7942 19564 7958
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 17696 7410 17724 7822
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18984 7546 19012 7754
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 19076 7478 19104 7822
rect 19708 7812 19760 7818
rect 19628 7772 19708 7800
rect 19214 7644 19522 7653
rect 19214 7642 19220 7644
rect 19276 7642 19300 7644
rect 19356 7642 19380 7644
rect 19436 7642 19460 7644
rect 19516 7642 19522 7644
rect 19276 7590 19278 7642
rect 19458 7590 19460 7642
rect 19214 7588 19220 7590
rect 19276 7588 19300 7590
rect 19356 7588 19380 7590
rect 19436 7588 19460 7590
rect 19516 7588 19522 7590
rect 19214 7579 19522 7588
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17696 6798 17724 7346
rect 19076 7002 19104 7414
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 17696 6322 17724 6734
rect 19628 6730 19656 7772
rect 19708 7754 19760 7760
rect 19996 7750 20024 8026
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19996 7546 20024 7686
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19214 6556 19522 6565
rect 19214 6554 19220 6556
rect 19276 6554 19300 6556
rect 19356 6554 19380 6556
rect 19436 6554 19460 6556
rect 19516 6554 19522 6556
rect 19276 6502 19278 6554
rect 19458 6502 19460 6554
rect 19214 6500 19220 6502
rect 19276 6500 19300 6502
rect 19356 6500 19380 6502
rect 19436 6500 19460 6502
rect 19516 6500 19522 6502
rect 19214 6491 19522 6500
rect 19628 6458 19656 6666
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17328 5914 17356 6258
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 19214 5468 19522 5477
rect 19214 5466 19220 5468
rect 19276 5466 19300 5468
rect 19356 5466 19380 5468
rect 19436 5466 19460 5468
rect 19516 5466 19522 5468
rect 19276 5414 19278 5466
rect 19458 5414 19460 5466
rect 19214 5412 19220 5414
rect 19276 5412 19300 5414
rect 19356 5412 19380 5414
rect 19436 5412 19460 5414
rect 19516 5412 19522 5414
rect 19214 5403 19522 5412
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14384 4214 14412 5306
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 16214 4924 16522 4933
rect 16214 4922 16220 4924
rect 16276 4922 16300 4924
rect 16356 4922 16380 4924
rect 16436 4922 16460 4924
rect 16516 4922 16522 4924
rect 16276 4870 16278 4922
rect 16458 4870 16460 4922
rect 16214 4868 16220 4870
rect 16276 4868 16300 4870
rect 16356 4868 16380 4870
rect 16436 4868 16460 4870
rect 16516 4868 16522 4870
rect 16214 4859 16522 4868
rect 20824 4865 20852 5170
rect 20810 4856 20866 4865
rect 20810 4791 20866 4800
rect 19214 4380 19522 4389
rect 19214 4378 19220 4380
rect 19276 4378 19300 4380
rect 19356 4378 19380 4380
rect 19436 4378 19460 4380
rect 19516 4378 19522 4380
rect 19276 4326 19278 4378
rect 19458 4326 19460 4378
rect 19214 4324 19220 4326
rect 19276 4324 19300 4326
rect 19356 4324 19380 4326
rect 19436 4324 19460 4326
rect 19516 4324 19522 4326
rect 19214 4315 19522 4324
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 14384 3466 14412 4150
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14372 3460 14424 3466
rect 14372 3402 14424 3408
rect 14752 3194 14780 3674
rect 14844 3602 14872 3878
rect 16214 3836 16522 3845
rect 16214 3834 16220 3836
rect 16276 3834 16300 3836
rect 16356 3834 16380 3836
rect 16436 3834 16460 3836
rect 16516 3834 16522 3836
rect 16276 3782 16278 3834
rect 16458 3782 16460 3834
rect 16214 3780 16220 3782
rect 16276 3780 16300 3782
rect 16356 3780 16380 3782
rect 16436 3780 16460 3782
rect 16516 3780 16522 3782
rect 16214 3771 16522 3780
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14844 3466 15240 3482
rect 14832 3460 15240 3466
rect 14884 3454 15240 3460
rect 14832 3402 14884 3408
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14384 2650 14412 2926
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 15212 2446 15240 3454
rect 19214 3292 19522 3301
rect 19214 3290 19220 3292
rect 19276 3290 19300 3292
rect 19356 3290 19380 3292
rect 19436 3290 19460 3292
rect 19516 3290 19522 3292
rect 19276 3238 19278 3290
rect 19458 3238 19460 3290
rect 19214 3236 19220 3238
rect 19276 3236 19300 3238
rect 19356 3236 19380 3238
rect 19436 3236 19460 3238
rect 19516 3236 19522 3238
rect 19214 3227 19522 3236
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 16214 2748 16522 2757
rect 16214 2746 16220 2748
rect 16276 2746 16300 2748
rect 16356 2746 16380 2748
rect 16436 2746 16460 2748
rect 16516 2746 16522 2748
rect 16276 2694 16278 2746
rect 16458 2694 16460 2746
rect 16214 2692 16220 2694
rect 16276 2692 16300 2694
rect 16356 2692 16380 2694
rect 16436 2692 16460 2694
rect 16516 2692 16522 2694
rect 16214 2683 16522 2692
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 13214 2204 13522 2213
rect 13214 2202 13220 2204
rect 13276 2202 13300 2204
rect 13356 2202 13380 2204
rect 13436 2202 13460 2204
rect 13516 2202 13522 2204
rect 13276 2150 13278 2202
rect 13458 2150 13460 2202
rect 13214 2148 13220 2150
rect 13276 2148 13300 2150
rect 13356 2148 13380 2150
rect 13436 2148 13460 2150
rect 13516 2148 13522 2150
rect 13214 2139 13522 2148
rect 15580 1170 15608 2314
rect 19214 2204 19522 2213
rect 19214 2202 19220 2204
rect 19276 2202 19300 2204
rect 19356 2202 19380 2204
rect 19436 2202 19460 2204
rect 19516 2202 19522 2204
rect 19276 2150 19278 2202
rect 19458 2150 19460 2202
rect 19214 2148 19220 2150
rect 19276 2148 19300 2150
rect 19356 2148 19380 2150
rect 19436 2148 19460 2150
rect 19516 2148 19522 2150
rect 19214 2139 19522 2148
rect 15488 1142 15608 1170
rect 15488 800 15516 1142
rect 20640 800 20668 2858
rect 10428 734 10640 762
rect 15474 0 15530 800
rect 20626 0 20682 800
<< via2 >>
rect 3606 21800 3662 21856
rect 938 16360 994 16416
rect 1398 10920 1454 10976
rect 1398 5480 1454 5536
rect 7220 21786 7276 21788
rect 7300 21786 7356 21788
rect 7380 21786 7436 21788
rect 7460 21786 7516 21788
rect 7220 21734 7266 21786
rect 7266 21734 7276 21786
rect 7300 21734 7330 21786
rect 7330 21734 7342 21786
rect 7342 21734 7356 21786
rect 7380 21734 7394 21786
rect 7394 21734 7406 21786
rect 7406 21734 7436 21786
rect 7460 21734 7470 21786
rect 7470 21734 7516 21786
rect 7220 21732 7276 21734
rect 7300 21732 7356 21734
rect 7380 21732 7436 21734
rect 7460 21732 7516 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 13220 21786 13276 21788
rect 13300 21786 13356 21788
rect 13380 21786 13436 21788
rect 13460 21786 13516 21788
rect 13220 21734 13266 21786
rect 13266 21734 13276 21786
rect 13300 21734 13330 21786
rect 13330 21734 13342 21786
rect 13342 21734 13356 21786
rect 13380 21734 13394 21786
rect 13394 21734 13406 21786
rect 13406 21734 13436 21786
rect 13460 21734 13470 21786
rect 13470 21734 13516 21786
rect 13220 21732 13276 21734
rect 13300 21732 13356 21734
rect 13380 21732 13436 21734
rect 13460 21732 13516 21734
rect 19220 21786 19276 21788
rect 19300 21786 19356 21788
rect 19380 21786 19436 21788
rect 19460 21786 19516 21788
rect 19220 21734 19266 21786
rect 19266 21734 19276 21786
rect 19300 21734 19330 21786
rect 19330 21734 19342 21786
rect 19342 21734 19356 21786
rect 19380 21734 19394 21786
rect 19394 21734 19406 21786
rect 19406 21734 19436 21786
rect 19460 21734 19470 21786
rect 19470 21734 19516 21786
rect 19220 21732 19276 21734
rect 19300 21732 19356 21734
rect 19380 21732 19436 21734
rect 19460 21732 19516 21734
rect 10220 21242 10276 21244
rect 10300 21242 10356 21244
rect 10380 21242 10436 21244
rect 10460 21242 10516 21244
rect 10220 21190 10266 21242
rect 10266 21190 10276 21242
rect 10300 21190 10330 21242
rect 10330 21190 10342 21242
rect 10342 21190 10356 21242
rect 10380 21190 10394 21242
rect 10394 21190 10406 21242
rect 10406 21190 10436 21242
rect 10460 21190 10470 21242
rect 10470 21190 10516 21242
rect 10220 21188 10276 21190
rect 10300 21188 10356 21190
rect 10380 21188 10436 21190
rect 10460 21188 10516 21190
rect 7220 20698 7276 20700
rect 7300 20698 7356 20700
rect 7380 20698 7436 20700
rect 7460 20698 7516 20700
rect 7220 20646 7266 20698
rect 7266 20646 7276 20698
rect 7300 20646 7330 20698
rect 7330 20646 7342 20698
rect 7342 20646 7356 20698
rect 7380 20646 7394 20698
rect 7394 20646 7406 20698
rect 7406 20646 7436 20698
rect 7460 20646 7470 20698
rect 7470 20646 7516 20698
rect 7220 20644 7276 20646
rect 7300 20644 7356 20646
rect 7380 20644 7436 20646
rect 7460 20644 7516 20646
rect 7220 19610 7276 19612
rect 7300 19610 7356 19612
rect 7380 19610 7436 19612
rect 7460 19610 7516 19612
rect 7220 19558 7266 19610
rect 7266 19558 7276 19610
rect 7300 19558 7330 19610
rect 7330 19558 7342 19610
rect 7342 19558 7356 19610
rect 7380 19558 7394 19610
rect 7394 19558 7406 19610
rect 7406 19558 7436 19610
rect 7460 19558 7470 19610
rect 7470 19558 7516 19610
rect 7220 19556 7276 19558
rect 7300 19556 7356 19558
rect 7380 19556 7436 19558
rect 7460 19556 7516 19558
rect 7220 18522 7276 18524
rect 7300 18522 7356 18524
rect 7380 18522 7436 18524
rect 7460 18522 7516 18524
rect 7220 18470 7266 18522
rect 7266 18470 7276 18522
rect 7300 18470 7330 18522
rect 7330 18470 7342 18522
rect 7342 18470 7356 18522
rect 7380 18470 7394 18522
rect 7394 18470 7406 18522
rect 7406 18470 7436 18522
rect 7460 18470 7470 18522
rect 7470 18470 7516 18522
rect 7220 18468 7276 18470
rect 7300 18468 7356 18470
rect 7380 18468 7436 18470
rect 7460 18468 7516 18470
rect 7220 17434 7276 17436
rect 7300 17434 7356 17436
rect 7380 17434 7436 17436
rect 7460 17434 7516 17436
rect 7220 17382 7266 17434
rect 7266 17382 7276 17434
rect 7300 17382 7330 17434
rect 7330 17382 7342 17434
rect 7342 17382 7356 17434
rect 7380 17382 7394 17434
rect 7394 17382 7406 17434
rect 7406 17382 7436 17434
rect 7460 17382 7470 17434
rect 7470 17382 7516 17434
rect 7220 17380 7276 17382
rect 7300 17380 7356 17382
rect 7380 17380 7436 17382
rect 7460 17380 7516 17382
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 7220 16346 7276 16348
rect 7300 16346 7356 16348
rect 7380 16346 7436 16348
rect 7460 16346 7516 16348
rect 7220 16294 7266 16346
rect 7266 16294 7276 16346
rect 7300 16294 7330 16346
rect 7330 16294 7342 16346
rect 7342 16294 7356 16346
rect 7380 16294 7394 16346
rect 7394 16294 7406 16346
rect 7406 16294 7436 16346
rect 7460 16294 7470 16346
rect 7470 16294 7516 16346
rect 7220 16292 7276 16294
rect 7300 16292 7356 16294
rect 7380 16292 7436 16294
rect 7460 16292 7516 16294
rect 7220 15258 7276 15260
rect 7300 15258 7356 15260
rect 7380 15258 7436 15260
rect 7460 15258 7516 15260
rect 7220 15206 7266 15258
rect 7266 15206 7276 15258
rect 7300 15206 7330 15258
rect 7330 15206 7342 15258
rect 7342 15206 7356 15258
rect 7380 15206 7394 15258
rect 7394 15206 7406 15258
rect 7406 15206 7436 15258
rect 7460 15206 7470 15258
rect 7470 15206 7516 15258
rect 7220 15204 7276 15206
rect 7300 15204 7356 15206
rect 7380 15204 7436 15206
rect 7460 15204 7516 15206
rect 7220 14170 7276 14172
rect 7300 14170 7356 14172
rect 7380 14170 7436 14172
rect 7460 14170 7516 14172
rect 7220 14118 7266 14170
rect 7266 14118 7276 14170
rect 7300 14118 7330 14170
rect 7330 14118 7342 14170
rect 7342 14118 7356 14170
rect 7380 14118 7394 14170
rect 7394 14118 7406 14170
rect 7406 14118 7436 14170
rect 7460 14118 7470 14170
rect 7470 14118 7516 14170
rect 7220 14116 7276 14118
rect 7300 14116 7356 14118
rect 7380 14116 7436 14118
rect 7460 14116 7516 14118
rect 7220 13082 7276 13084
rect 7300 13082 7356 13084
rect 7380 13082 7436 13084
rect 7460 13082 7516 13084
rect 7220 13030 7266 13082
rect 7266 13030 7276 13082
rect 7300 13030 7330 13082
rect 7330 13030 7342 13082
rect 7342 13030 7356 13082
rect 7380 13030 7394 13082
rect 7394 13030 7406 13082
rect 7406 13030 7436 13082
rect 7460 13030 7470 13082
rect 7470 13030 7516 13082
rect 7220 13028 7276 13030
rect 7300 13028 7356 13030
rect 7380 13028 7436 13030
rect 7460 13028 7516 13030
rect 7220 11994 7276 11996
rect 7300 11994 7356 11996
rect 7380 11994 7436 11996
rect 7460 11994 7516 11996
rect 7220 11942 7266 11994
rect 7266 11942 7276 11994
rect 7300 11942 7330 11994
rect 7330 11942 7342 11994
rect 7342 11942 7356 11994
rect 7380 11942 7394 11994
rect 7394 11942 7406 11994
rect 7406 11942 7436 11994
rect 7460 11942 7470 11994
rect 7470 11942 7516 11994
rect 7220 11940 7276 11942
rect 7300 11940 7356 11942
rect 7380 11940 7436 11942
rect 7460 11940 7516 11942
rect 7220 10906 7276 10908
rect 7300 10906 7356 10908
rect 7380 10906 7436 10908
rect 7460 10906 7516 10908
rect 7220 10854 7266 10906
rect 7266 10854 7276 10906
rect 7300 10854 7330 10906
rect 7330 10854 7342 10906
rect 7342 10854 7356 10906
rect 7380 10854 7394 10906
rect 7394 10854 7406 10906
rect 7406 10854 7436 10906
rect 7460 10854 7470 10906
rect 7470 10854 7516 10906
rect 7220 10852 7276 10854
rect 7300 10852 7356 10854
rect 7380 10852 7436 10854
rect 7460 10852 7516 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 7220 9818 7276 9820
rect 7300 9818 7356 9820
rect 7380 9818 7436 9820
rect 7460 9818 7516 9820
rect 7220 9766 7266 9818
rect 7266 9766 7276 9818
rect 7300 9766 7330 9818
rect 7330 9766 7342 9818
rect 7342 9766 7356 9818
rect 7380 9766 7394 9818
rect 7394 9766 7406 9818
rect 7406 9766 7436 9818
rect 7460 9766 7470 9818
rect 7470 9766 7516 9818
rect 7220 9764 7276 9766
rect 7300 9764 7356 9766
rect 7380 9764 7436 9766
rect 7460 9764 7516 9766
rect 7220 8730 7276 8732
rect 7300 8730 7356 8732
rect 7380 8730 7436 8732
rect 7460 8730 7516 8732
rect 7220 8678 7266 8730
rect 7266 8678 7276 8730
rect 7300 8678 7330 8730
rect 7330 8678 7342 8730
rect 7342 8678 7356 8730
rect 7380 8678 7394 8730
rect 7394 8678 7406 8730
rect 7406 8678 7436 8730
rect 7460 8678 7470 8730
rect 7470 8678 7516 8730
rect 7220 8676 7276 8678
rect 7300 8676 7356 8678
rect 7380 8676 7436 8678
rect 7460 8676 7516 8678
rect 7220 7642 7276 7644
rect 7300 7642 7356 7644
rect 7380 7642 7436 7644
rect 7460 7642 7516 7644
rect 7220 7590 7266 7642
rect 7266 7590 7276 7642
rect 7300 7590 7330 7642
rect 7330 7590 7342 7642
rect 7342 7590 7356 7642
rect 7380 7590 7394 7642
rect 7394 7590 7406 7642
rect 7406 7590 7436 7642
rect 7460 7590 7470 7642
rect 7470 7590 7516 7642
rect 7220 7588 7276 7590
rect 7300 7588 7356 7590
rect 7380 7588 7436 7590
rect 7460 7588 7516 7590
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 7220 6554 7276 6556
rect 7300 6554 7356 6556
rect 7380 6554 7436 6556
rect 7460 6554 7516 6556
rect 7220 6502 7266 6554
rect 7266 6502 7276 6554
rect 7300 6502 7330 6554
rect 7330 6502 7342 6554
rect 7342 6502 7356 6554
rect 7380 6502 7394 6554
rect 7394 6502 7406 6554
rect 7406 6502 7436 6554
rect 7460 6502 7470 6554
rect 7470 6502 7516 6554
rect 7220 6500 7276 6502
rect 7300 6500 7356 6502
rect 7380 6500 7436 6502
rect 7460 6500 7516 6502
rect 10220 20154 10276 20156
rect 10300 20154 10356 20156
rect 10380 20154 10436 20156
rect 10460 20154 10516 20156
rect 10220 20102 10266 20154
rect 10266 20102 10276 20154
rect 10300 20102 10330 20154
rect 10330 20102 10342 20154
rect 10342 20102 10356 20154
rect 10380 20102 10394 20154
rect 10394 20102 10406 20154
rect 10406 20102 10436 20154
rect 10460 20102 10470 20154
rect 10470 20102 10516 20154
rect 10220 20100 10276 20102
rect 10300 20100 10356 20102
rect 10380 20100 10436 20102
rect 10460 20100 10516 20102
rect 10220 19066 10276 19068
rect 10300 19066 10356 19068
rect 10380 19066 10436 19068
rect 10460 19066 10516 19068
rect 10220 19014 10266 19066
rect 10266 19014 10276 19066
rect 10300 19014 10330 19066
rect 10330 19014 10342 19066
rect 10342 19014 10356 19066
rect 10380 19014 10394 19066
rect 10394 19014 10406 19066
rect 10406 19014 10436 19066
rect 10460 19014 10470 19066
rect 10470 19014 10516 19066
rect 10220 19012 10276 19014
rect 10300 19012 10356 19014
rect 10380 19012 10436 19014
rect 10460 19012 10516 19014
rect 13220 20698 13276 20700
rect 13300 20698 13356 20700
rect 13380 20698 13436 20700
rect 13460 20698 13516 20700
rect 13220 20646 13266 20698
rect 13266 20646 13276 20698
rect 13300 20646 13330 20698
rect 13330 20646 13342 20698
rect 13342 20646 13356 20698
rect 13380 20646 13394 20698
rect 13394 20646 13406 20698
rect 13406 20646 13436 20698
rect 13460 20646 13470 20698
rect 13470 20646 13516 20698
rect 13220 20644 13276 20646
rect 13300 20644 13356 20646
rect 13380 20644 13436 20646
rect 13460 20644 13516 20646
rect 16220 21242 16276 21244
rect 16300 21242 16356 21244
rect 16380 21242 16436 21244
rect 16460 21242 16516 21244
rect 16220 21190 16266 21242
rect 16266 21190 16276 21242
rect 16300 21190 16330 21242
rect 16330 21190 16342 21242
rect 16342 21190 16356 21242
rect 16380 21190 16394 21242
rect 16394 21190 16406 21242
rect 16406 21190 16436 21242
rect 16460 21190 16470 21242
rect 16470 21190 16516 21242
rect 16220 21188 16276 21190
rect 16300 21188 16356 21190
rect 16380 21188 16436 21190
rect 16460 21188 16516 21190
rect 13220 19610 13276 19612
rect 13300 19610 13356 19612
rect 13380 19610 13436 19612
rect 13460 19610 13516 19612
rect 13220 19558 13266 19610
rect 13266 19558 13276 19610
rect 13300 19558 13330 19610
rect 13330 19558 13342 19610
rect 13342 19558 13356 19610
rect 13380 19558 13394 19610
rect 13394 19558 13406 19610
rect 13406 19558 13436 19610
rect 13460 19558 13470 19610
rect 13470 19558 13516 19610
rect 13220 19556 13276 19558
rect 13300 19556 13356 19558
rect 13380 19556 13436 19558
rect 13460 19556 13516 19558
rect 10220 17978 10276 17980
rect 10300 17978 10356 17980
rect 10380 17978 10436 17980
rect 10460 17978 10516 17980
rect 10220 17926 10266 17978
rect 10266 17926 10276 17978
rect 10300 17926 10330 17978
rect 10330 17926 10342 17978
rect 10342 17926 10356 17978
rect 10380 17926 10394 17978
rect 10394 17926 10406 17978
rect 10406 17926 10436 17978
rect 10460 17926 10470 17978
rect 10470 17926 10516 17978
rect 10220 17924 10276 17926
rect 10300 17924 10356 17926
rect 10380 17924 10436 17926
rect 10460 17924 10516 17926
rect 10220 16890 10276 16892
rect 10300 16890 10356 16892
rect 10380 16890 10436 16892
rect 10460 16890 10516 16892
rect 10220 16838 10266 16890
rect 10266 16838 10276 16890
rect 10300 16838 10330 16890
rect 10330 16838 10342 16890
rect 10342 16838 10356 16890
rect 10380 16838 10394 16890
rect 10394 16838 10406 16890
rect 10406 16838 10436 16890
rect 10460 16838 10470 16890
rect 10470 16838 10516 16890
rect 10220 16836 10276 16838
rect 10300 16836 10356 16838
rect 10380 16836 10436 16838
rect 10460 16836 10516 16838
rect 10220 15802 10276 15804
rect 10300 15802 10356 15804
rect 10380 15802 10436 15804
rect 10460 15802 10516 15804
rect 10220 15750 10266 15802
rect 10266 15750 10276 15802
rect 10300 15750 10330 15802
rect 10330 15750 10342 15802
rect 10342 15750 10356 15802
rect 10380 15750 10394 15802
rect 10394 15750 10406 15802
rect 10406 15750 10436 15802
rect 10460 15750 10470 15802
rect 10470 15750 10516 15802
rect 10220 15748 10276 15750
rect 10300 15748 10356 15750
rect 10380 15748 10436 15750
rect 10460 15748 10516 15750
rect 13220 18522 13276 18524
rect 13300 18522 13356 18524
rect 13380 18522 13436 18524
rect 13460 18522 13516 18524
rect 13220 18470 13266 18522
rect 13266 18470 13276 18522
rect 13300 18470 13330 18522
rect 13330 18470 13342 18522
rect 13342 18470 13356 18522
rect 13380 18470 13394 18522
rect 13394 18470 13406 18522
rect 13406 18470 13436 18522
rect 13460 18470 13470 18522
rect 13470 18470 13516 18522
rect 13220 18468 13276 18470
rect 13300 18468 13356 18470
rect 13380 18468 13436 18470
rect 13460 18468 13516 18470
rect 13220 17434 13276 17436
rect 13300 17434 13356 17436
rect 13380 17434 13436 17436
rect 13460 17434 13516 17436
rect 13220 17382 13266 17434
rect 13266 17382 13276 17434
rect 13300 17382 13330 17434
rect 13330 17382 13342 17434
rect 13342 17382 13356 17434
rect 13380 17382 13394 17434
rect 13394 17382 13406 17434
rect 13406 17382 13436 17434
rect 13460 17382 13470 17434
rect 13470 17382 13516 17434
rect 13220 17380 13276 17382
rect 13300 17380 13356 17382
rect 13380 17380 13436 17382
rect 13460 17380 13516 17382
rect 10220 14714 10276 14716
rect 10300 14714 10356 14716
rect 10380 14714 10436 14716
rect 10460 14714 10516 14716
rect 10220 14662 10266 14714
rect 10266 14662 10276 14714
rect 10300 14662 10330 14714
rect 10330 14662 10342 14714
rect 10342 14662 10356 14714
rect 10380 14662 10394 14714
rect 10394 14662 10406 14714
rect 10406 14662 10436 14714
rect 10460 14662 10470 14714
rect 10470 14662 10516 14714
rect 10220 14660 10276 14662
rect 10300 14660 10356 14662
rect 10380 14660 10436 14662
rect 10460 14660 10516 14662
rect 10220 13626 10276 13628
rect 10300 13626 10356 13628
rect 10380 13626 10436 13628
rect 10460 13626 10516 13628
rect 10220 13574 10266 13626
rect 10266 13574 10276 13626
rect 10300 13574 10330 13626
rect 10330 13574 10342 13626
rect 10342 13574 10356 13626
rect 10380 13574 10394 13626
rect 10394 13574 10406 13626
rect 10406 13574 10436 13626
rect 10460 13574 10470 13626
rect 10470 13574 10516 13626
rect 10220 13572 10276 13574
rect 10300 13572 10356 13574
rect 10380 13572 10436 13574
rect 10460 13572 10516 13574
rect 13220 16346 13276 16348
rect 13300 16346 13356 16348
rect 13380 16346 13436 16348
rect 13460 16346 13516 16348
rect 13220 16294 13266 16346
rect 13266 16294 13276 16346
rect 13300 16294 13330 16346
rect 13330 16294 13342 16346
rect 13342 16294 13356 16346
rect 13380 16294 13394 16346
rect 13394 16294 13406 16346
rect 13406 16294 13436 16346
rect 13460 16294 13470 16346
rect 13470 16294 13516 16346
rect 13220 16292 13276 16294
rect 13300 16292 13356 16294
rect 13380 16292 13436 16294
rect 13460 16292 13516 16294
rect 13220 15258 13276 15260
rect 13300 15258 13356 15260
rect 13380 15258 13436 15260
rect 13460 15258 13516 15260
rect 13220 15206 13266 15258
rect 13266 15206 13276 15258
rect 13300 15206 13330 15258
rect 13330 15206 13342 15258
rect 13342 15206 13356 15258
rect 13380 15206 13394 15258
rect 13394 15206 13406 15258
rect 13406 15206 13436 15258
rect 13460 15206 13470 15258
rect 13470 15206 13516 15258
rect 13220 15204 13276 15206
rect 13300 15204 13356 15206
rect 13380 15204 13436 15206
rect 13460 15204 13516 15206
rect 13220 14170 13276 14172
rect 13300 14170 13356 14172
rect 13380 14170 13436 14172
rect 13460 14170 13516 14172
rect 13220 14118 13266 14170
rect 13266 14118 13276 14170
rect 13300 14118 13330 14170
rect 13330 14118 13342 14170
rect 13342 14118 13356 14170
rect 13380 14118 13394 14170
rect 13394 14118 13406 14170
rect 13406 14118 13436 14170
rect 13460 14118 13470 14170
rect 13470 14118 13516 14170
rect 13220 14116 13276 14118
rect 13300 14116 13356 14118
rect 13380 14116 13436 14118
rect 13460 14116 13516 14118
rect 16220 20154 16276 20156
rect 16300 20154 16356 20156
rect 16380 20154 16436 20156
rect 16460 20154 16516 20156
rect 16220 20102 16266 20154
rect 16266 20102 16276 20154
rect 16300 20102 16330 20154
rect 16330 20102 16342 20154
rect 16342 20102 16356 20154
rect 16380 20102 16394 20154
rect 16394 20102 16406 20154
rect 16406 20102 16436 20154
rect 16460 20102 16470 20154
rect 16470 20102 16516 20154
rect 16220 20100 16276 20102
rect 16300 20100 16356 20102
rect 16380 20100 16436 20102
rect 16460 20100 16516 20102
rect 16220 19066 16276 19068
rect 16300 19066 16356 19068
rect 16380 19066 16436 19068
rect 16460 19066 16516 19068
rect 16220 19014 16266 19066
rect 16266 19014 16276 19066
rect 16300 19014 16330 19066
rect 16330 19014 16342 19066
rect 16342 19014 16356 19066
rect 16380 19014 16394 19066
rect 16394 19014 16406 19066
rect 16406 19014 16436 19066
rect 16460 19014 16470 19066
rect 16470 19014 16516 19066
rect 16220 19012 16276 19014
rect 16300 19012 16356 19014
rect 16380 19012 16436 19014
rect 16460 19012 16516 19014
rect 16220 17978 16276 17980
rect 16300 17978 16356 17980
rect 16380 17978 16436 17980
rect 16460 17978 16516 17980
rect 16220 17926 16266 17978
rect 16266 17926 16276 17978
rect 16300 17926 16330 17978
rect 16330 17926 16342 17978
rect 16342 17926 16356 17978
rect 16380 17926 16394 17978
rect 16394 17926 16406 17978
rect 16406 17926 16436 17978
rect 16460 17926 16470 17978
rect 16470 17926 16516 17978
rect 16220 17924 16276 17926
rect 16300 17924 16356 17926
rect 16380 17924 16436 17926
rect 16460 17924 16516 17926
rect 16220 16890 16276 16892
rect 16300 16890 16356 16892
rect 16380 16890 16436 16892
rect 16460 16890 16516 16892
rect 16220 16838 16266 16890
rect 16266 16838 16276 16890
rect 16300 16838 16330 16890
rect 16330 16838 16342 16890
rect 16342 16838 16356 16890
rect 16380 16838 16394 16890
rect 16394 16838 16406 16890
rect 16406 16838 16436 16890
rect 16460 16838 16470 16890
rect 16470 16838 16516 16890
rect 16220 16836 16276 16838
rect 16300 16836 16356 16838
rect 16380 16836 16436 16838
rect 16460 16836 16516 16838
rect 16220 15802 16276 15804
rect 16300 15802 16356 15804
rect 16380 15802 16436 15804
rect 16460 15802 16516 15804
rect 16220 15750 16266 15802
rect 16266 15750 16276 15802
rect 16300 15750 16330 15802
rect 16330 15750 16342 15802
rect 16342 15750 16356 15802
rect 16380 15750 16394 15802
rect 16394 15750 16406 15802
rect 16406 15750 16436 15802
rect 16460 15750 16470 15802
rect 16470 15750 16516 15802
rect 16220 15748 16276 15750
rect 16300 15748 16356 15750
rect 16380 15748 16436 15750
rect 16460 15748 16516 15750
rect 16220 14714 16276 14716
rect 16300 14714 16356 14716
rect 16380 14714 16436 14716
rect 16460 14714 16516 14716
rect 16220 14662 16266 14714
rect 16266 14662 16276 14714
rect 16300 14662 16330 14714
rect 16330 14662 16342 14714
rect 16342 14662 16356 14714
rect 16380 14662 16394 14714
rect 16394 14662 16406 14714
rect 16406 14662 16436 14714
rect 16460 14662 16470 14714
rect 16470 14662 16516 14714
rect 16220 14660 16276 14662
rect 16300 14660 16356 14662
rect 16380 14660 16436 14662
rect 16460 14660 16516 14662
rect 17038 15680 17094 15736
rect 10220 12538 10276 12540
rect 10300 12538 10356 12540
rect 10380 12538 10436 12540
rect 10460 12538 10516 12540
rect 10220 12486 10266 12538
rect 10266 12486 10276 12538
rect 10300 12486 10330 12538
rect 10330 12486 10342 12538
rect 10342 12486 10356 12538
rect 10380 12486 10394 12538
rect 10394 12486 10406 12538
rect 10406 12486 10436 12538
rect 10460 12486 10470 12538
rect 10470 12486 10516 12538
rect 10220 12484 10276 12486
rect 10300 12484 10356 12486
rect 10380 12484 10436 12486
rect 10460 12484 10516 12486
rect 10220 11450 10276 11452
rect 10300 11450 10356 11452
rect 10380 11450 10436 11452
rect 10460 11450 10516 11452
rect 10220 11398 10266 11450
rect 10266 11398 10276 11450
rect 10300 11398 10330 11450
rect 10330 11398 10342 11450
rect 10342 11398 10356 11450
rect 10380 11398 10394 11450
rect 10394 11398 10406 11450
rect 10406 11398 10436 11450
rect 10460 11398 10470 11450
rect 10470 11398 10516 11450
rect 10220 11396 10276 11398
rect 10300 11396 10356 11398
rect 10380 11396 10436 11398
rect 10460 11396 10516 11398
rect 7220 5466 7276 5468
rect 7300 5466 7356 5468
rect 7380 5466 7436 5468
rect 7460 5466 7516 5468
rect 7220 5414 7266 5466
rect 7266 5414 7276 5466
rect 7300 5414 7330 5466
rect 7330 5414 7342 5466
rect 7342 5414 7356 5466
rect 7380 5414 7394 5466
rect 7394 5414 7406 5466
rect 7406 5414 7436 5466
rect 7460 5414 7470 5466
rect 7470 5414 7516 5466
rect 7220 5412 7276 5414
rect 7300 5412 7356 5414
rect 7380 5412 7436 5414
rect 7460 5412 7516 5414
rect 7220 4378 7276 4380
rect 7300 4378 7356 4380
rect 7380 4378 7436 4380
rect 7460 4378 7516 4380
rect 7220 4326 7266 4378
rect 7266 4326 7276 4378
rect 7300 4326 7330 4378
rect 7330 4326 7342 4378
rect 7342 4326 7356 4378
rect 7380 4326 7394 4378
rect 7394 4326 7406 4378
rect 7406 4326 7436 4378
rect 7460 4326 7470 4378
rect 7470 4326 7516 4378
rect 7220 4324 7276 4326
rect 7300 4324 7356 4326
rect 7380 4324 7436 4326
rect 7460 4324 7516 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 7220 3290 7276 3292
rect 7300 3290 7356 3292
rect 7380 3290 7436 3292
rect 7460 3290 7516 3292
rect 7220 3238 7266 3290
rect 7266 3238 7276 3290
rect 7300 3238 7330 3290
rect 7330 3238 7342 3290
rect 7342 3238 7356 3290
rect 7380 3238 7394 3290
rect 7394 3238 7406 3290
rect 7406 3238 7436 3290
rect 7460 3238 7470 3290
rect 7470 3238 7516 3290
rect 7220 3236 7276 3238
rect 7300 3236 7356 3238
rect 7380 3236 7436 3238
rect 7460 3236 7516 3238
rect 10220 10362 10276 10364
rect 10300 10362 10356 10364
rect 10380 10362 10436 10364
rect 10460 10362 10516 10364
rect 10220 10310 10266 10362
rect 10266 10310 10276 10362
rect 10300 10310 10330 10362
rect 10330 10310 10342 10362
rect 10342 10310 10356 10362
rect 10380 10310 10394 10362
rect 10394 10310 10406 10362
rect 10406 10310 10436 10362
rect 10460 10310 10470 10362
rect 10470 10310 10516 10362
rect 10220 10308 10276 10310
rect 10300 10308 10356 10310
rect 10380 10308 10436 10310
rect 10460 10308 10516 10310
rect 10220 9274 10276 9276
rect 10300 9274 10356 9276
rect 10380 9274 10436 9276
rect 10460 9274 10516 9276
rect 10220 9222 10266 9274
rect 10266 9222 10276 9274
rect 10300 9222 10330 9274
rect 10330 9222 10342 9274
rect 10342 9222 10356 9274
rect 10380 9222 10394 9274
rect 10394 9222 10406 9274
rect 10406 9222 10436 9274
rect 10460 9222 10470 9274
rect 10470 9222 10516 9274
rect 10220 9220 10276 9222
rect 10300 9220 10356 9222
rect 10380 9220 10436 9222
rect 10460 9220 10516 9222
rect 10220 8186 10276 8188
rect 10300 8186 10356 8188
rect 10380 8186 10436 8188
rect 10460 8186 10516 8188
rect 10220 8134 10266 8186
rect 10266 8134 10276 8186
rect 10300 8134 10330 8186
rect 10330 8134 10342 8186
rect 10342 8134 10356 8186
rect 10380 8134 10394 8186
rect 10394 8134 10406 8186
rect 10406 8134 10436 8186
rect 10460 8134 10470 8186
rect 10470 8134 10516 8186
rect 10220 8132 10276 8134
rect 10300 8132 10356 8134
rect 10380 8132 10436 8134
rect 10460 8132 10516 8134
rect 13220 13082 13276 13084
rect 13300 13082 13356 13084
rect 13380 13082 13436 13084
rect 13460 13082 13516 13084
rect 13220 13030 13266 13082
rect 13266 13030 13276 13082
rect 13300 13030 13330 13082
rect 13330 13030 13342 13082
rect 13342 13030 13356 13082
rect 13380 13030 13394 13082
rect 13394 13030 13406 13082
rect 13406 13030 13436 13082
rect 13460 13030 13470 13082
rect 13470 13030 13516 13082
rect 13220 13028 13276 13030
rect 13300 13028 13356 13030
rect 13380 13028 13436 13030
rect 13460 13028 13516 13030
rect 13220 11994 13276 11996
rect 13300 11994 13356 11996
rect 13380 11994 13436 11996
rect 13460 11994 13516 11996
rect 13220 11942 13266 11994
rect 13266 11942 13276 11994
rect 13300 11942 13330 11994
rect 13330 11942 13342 11994
rect 13342 11942 13356 11994
rect 13380 11942 13394 11994
rect 13394 11942 13406 11994
rect 13406 11942 13436 11994
rect 13460 11942 13470 11994
rect 13470 11942 13516 11994
rect 13220 11940 13276 11942
rect 13300 11940 13356 11942
rect 13380 11940 13436 11942
rect 13460 11940 13516 11942
rect 16220 13626 16276 13628
rect 16300 13626 16356 13628
rect 16380 13626 16436 13628
rect 16460 13626 16516 13628
rect 16220 13574 16266 13626
rect 16266 13574 16276 13626
rect 16300 13574 16330 13626
rect 16330 13574 16342 13626
rect 16342 13574 16356 13626
rect 16380 13574 16394 13626
rect 16394 13574 16406 13626
rect 16406 13574 16436 13626
rect 16460 13574 16470 13626
rect 16470 13574 16516 13626
rect 16220 13572 16276 13574
rect 16300 13572 16356 13574
rect 16380 13572 16436 13574
rect 16460 13572 16516 13574
rect 16220 12538 16276 12540
rect 16300 12538 16356 12540
rect 16380 12538 16436 12540
rect 16460 12538 16516 12540
rect 16220 12486 16266 12538
rect 16266 12486 16276 12538
rect 16300 12486 16330 12538
rect 16330 12486 16342 12538
rect 16342 12486 16356 12538
rect 16380 12486 16394 12538
rect 16394 12486 16406 12538
rect 16406 12486 16436 12538
rect 16460 12486 16470 12538
rect 16470 12486 16516 12538
rect 16220 12484 16276 12486
rect 16300 12484 16356 12486
rect 16380 12484 16436 12486
rect 16460 12484 16516 12486
rect 13220 10906 13276 10908
rect 13300 10906 13356 10908
rect 13380 10906 13436 10908
rect 13460 10906 13516 10908
rect 13220 10854 13266 10906
rect 13266 10854 13276 10906
rect 13300 10854 13330 10906
rect 13330 10854 13342 10906
rect 13342 10854 13356 10906
rect 13380 10854 13394 10906
rect 13394 10854 13406 10906
rect 13406 10854 13436 10906
rect 13460 10854 13470 10906
rect 13470 10854 13516 10906
rect 13220 10852 13276 10854
rect 13300 10852 13356 10854
rect 13380 10852 13436 10854
rect 13460 10852 13516 10854
rect 10220 7098 10276 7100
rect 10300 7098 10356 7100
rect 10380 7098 10436 7100
rect 10460 7098 10516 7100
rect 10220 7046 10266 7098
rect 10266 7046 10276 7098
rect 10300 7046 10330 7098
rect 10330 7046 10342 7098
rect 10342 7046 10356 7098
rect 10380 7046 10394 7098
rect 10394 7046 10406 7098
rect 10406 7046 10436 7098
rect 10460 7046 10470 7098
rect 10470 7046 10516 7098
rect 10220 7044 10276 7046
rect 10300 7044 10356 7046
rect 10380 7044 10436 7046
rect 10460 7044 10516 7046
rect 10220 6010 10276 6012
rect 10300 6010 10356 6012
rect 10380 6010 10436 6012
rect 10460 6010 10516 6012
rect 10220 5958 10266 6010
rect 10266 5958 10276 6010
rect 10300 5958 10330 6010
rect 10330 5958 10342 6010
rect 10342 5958 10356 6010
rect 10380 5958 10394 6010
rect 10394 5958 10406 6010
rect 10406 5958 10436 6010
rect 10460 5958 10470 6010
rect 10470 5958 10516 6010
rect 10220 5956 10276 5958
rect 10300 5956 10356 5958
rect 10380 5956 10436 5958
rect 10460 5956 10516 5958
rect 10220 4922 10276 4924
rect 10300 4922 10356 4924
rect 10380 4922 10436 4924
rect 10460 4922 10516 4924
rect 10220 4870 10266 4922
rect 10266 4870 10276 4922
rect 10300 4870 10330 4922
rect 10330 4870 10342 4922
rect 10342 4870 10356 4922
rect 10380 4870 10394 4922
rect 10394 4870 10406 4922
rect 10406 4870 10436 4922
rect 10460 4870 10470 4922
rect 10470 4870 10516 4922
rect 10220 4868 10276 4870
rect 10300 4868 10356 4870
rect 10380 4868 10436 4870
rect 10460 4868 10516 4870
rect 10220 3834 10276 3836
rect 10300 3834 10356 3836
rect 10380 3834 10436 3836
rect 10460 3834 10516 3836
rect 10220 3782 10266 3834
rect 10266 3782 10276 3834
rect 10300 3782 10330 3834
rect 10330 3782 10342 3834
rect 10342 3782 10356 3834
rect 10380 3782 10394 3834
rect 10394 3782 10406 3834
rect 10406 3782 10436 3834
rect 10460 3782 10470 3834
rect 10470 3782 10516 3834
rect 10220 3780 10276 3782
rect 10300 3780 10356 3782
rect 10380 3780 10436 3782
rect 10460 3780 10516 3782
rect 10220 2746 10276 2748
rect 10300 2746 10356 2748
rect 10380 2746 10436 2748
rect 10460 2746 10516 2748
rect 10220 2694 10266 2746
rect 10266 2694 10276 2746
rect 10300 2694 10330 2746
rect 10330 2694 10342 2746
rect 10342 2694 10356 2746
rect 10380 2694 10394 2746
rect 10394 2694 10406 2746
rect 10406 2694 10436 2746
rect 10460 2694 10470 2746
rect 10470 2694 10516 2746
rect 10220 2692 10276 2694
rect 10300 2692 10356 2694
rect 10380 2692 10436 2694
rect 10460 2692 10516 2694
rect 7220 2202 7276 2204
rect 7300 2202 7356 2204
rect 7380 2202 7436 2204
rect 7460 2202 7516 2204
rect 7220 2150 7266 2202
rect 7266 2150 7276 2202
rect 7300 2150 7330 2202
rect 7330 2150 7342 2202
rect 7342 2150 7356 2202
rect 7380 2150 7394 2202
rect 7394 2150 7406 2202
rect 7406 2150 7436 2202
rect 7460 2150 7470 2202
rect 7470 2150 7516 2202
rect 7220 2148 7276 2150
rect 7300 2148 7356 2150
rect 7380 2148 7436 2150
rect 7460 2148 7516 2150
rect 13220 9818 13276 9820
rect 13300 9818 13356 9820
rect 13380 9818 13436 9820
rect 13460 9818 13516 9820
rect 13220 9766 13266 9818
rect 13266 9766 13276 9818
rect 13300 9766 13330 9818
rect 13330 9766 13342 9818
rect 13342 9766 13356 9818
rect 13380 9766 13394 9818
rect 13394 9766 13406 9818
rect 13406 9766 13436 9818
rect 13460 9766 13470 9818
rect 13470 9766 13516 9818
rect 13220 9764 13276 9766
rect 13300 9764 13356 9766
rect 13380 9764 13436 9766
rect 13460 9764 13516 9766
rect 13220 8730 13276 8732
rect 13300 8730 13356 8732
rect 13380 8730 13436 8732
rect 13460 8730 13516 8732
rect 13220 8678 13266 8730
rect 13266 8678 13276 8730
rect 13300 8678 13330 8730
rect 13330 8678 13342 8730
rect 13342 8678 13356 8730
rect 13380 8678 13394 8730
rect 13394 8678 13406 8730
rect 13406 8678 13436 8730
rect 13460 8678 13470 8730
rect 13470 8678 13516 8730
rect 13220 8676 13276 8678
rect 13300 8676 13356 8678
rect 13380 8676 13436 8678
rect 13460 8676 13516 8678
rect 13220 7642 13276 7644
rect 13300 7642 13356 7644
rect 13380 7642 13436 7644
rect 13460 7642 13516 7644
rect 13220 7590 13266 7642
rect 13266 7590 13276 7642
rect 13300 7590 13330 7642
rect 13330 7590 13342 7642
rect 13342 7590 13356 7642
rect 13380 7590 13394 7642
rect 13394 7590 13406 7642
rect 13406 7590 13436 7642
rect 13460 7590 13470 7642
rect 13470 7590 13516 7642
rect 13220 7588 13276 7590
rect 13300 7588 13356 7590
rect 13380 7588 13436 7590
rect 13460 7588 13516 7590
rect 13220 6554 13276 6556
rect 13300 6554 13356 6556
rect 13380 6554 13436 6556
rect 13460 6554 13516 6556
rect 13220 6502 13266 6554
rect 13266 6502 13276 6554
rect 13300 6502 13330 6554
rect 13330 6502 13342 6554
rect 13342 6502 13356 6554
rect 13380 6502 13394 6554
rect 13394 6502 13406 6554
rect 13406 6502 13436 6554
rect 13460 6502 13470 6554
rect 13470 6502 13516 6554
rect 13220 6500 13276 6502
rect 13300 6500 13356 6502
rect 13380 6500 13436 6502
rect 13460 6500 13516 6502
rect 13220 5466 13276 5468
rect 13300 5466 13356 5468
rect 13380 5466 13436 5468
rect 13460 5466 13516 5468
rect 13220 5414 13266 5466
rect 13266 5414 13276 5466
rect 13300 5414 13330 5466
rect 13330 5414 13342 5466
rect 13342 5414 13356 5466
rect 13380 5414 13394 5466
rect 13394 5414 13406 5466
rect 13406 5414 13436 5466
rect 13460 5414 13470 5466
rect 13470 5414 13516 5466
rect 13220 5412 13276 5414
rect 13300 5412 13356 5414
rect 13380 5412 13436 5414
rect 13460 5412 13516 5414
rect 16220 11450 16276 11452
rect 16300 11450 16356 11452
rect 16380 11450 16436 11452
rect 16460 11450 16516 11452
rect 16220 11398 16266 11450
rect 16266 11398 16276 11450
rect 16300 11398 16330 11450
rect 16330 11398 16342 11450
rect 16342 11398 16356 11450
rect 16380 11398 16394 11450
rect 16394 11398 16406 11450
rect 16406 11398 16436 11450
rect 16460 11398 16470 11450
rect 16470 11398 16516 11450
rect 16220 11396 16276 11398
rect 16300 11396 16356 11398
rect 16380 11396 16436 11398
rect 16460 11396 16516 11398
rect 19220 20698 19276 20700
rect 19300 20698 19356 20700
rect 19380 20698 19436 20700
rect 19460 20698 19516 20700
rect 19220 20646 19266 20698
rect 19266 20646 19276 20698
rect 19300 20646 19330 20698
rect 19330 20646 19342 20698
rect 19342 20646 19356 20698
rect 19380 20646 19394 20698
rect 19394 20646 19406 20698
rect 19406 20646 19436 20698
rect 19460 20646 19470 20698
rect 19470 20646 19516 20698
rect 19220 20644 19276 20646
rect 19300 20644 19356 20646
rect 19380 20644 19436 20646
rect 19460 20644 19516 20646
rect 19220 19610 19276 19612
rect 19300 19610 19356 19612
rect 19380 19610 19436 19612
rect 19460 19610 19516 19612
rect 19220 19558 19266 19610
rect 19266 19558 19276 19610
rect 19300 19558 19330 19610
rect 19330 19558 19342 19610
rect 19342 19558 19356 19610
rect 19380 19558 19394 19610
rect 19394 19558 19406 19610
rect 19406 19558 19436 19610
rect 19460 19558 19470 19610
rect 19470 19558 19516 19610
rect 19220 19556 19276 19558
rect 19300 19556 19356 19558
rect 19380 19556 19436 19558
rect 19460 19556 19516 19558
rect 19220 18522 19276 18524
rect 19300 18522 19356 18524
rect 19380 18522 19436 18524
rect 19460 18522 19516 18524
rect 19220 18470 19266 18522
rect 19266 18470 19276 18522
rect 19300 18470 19330 18522
rect 19330 18470 19342 18522
rect 19342 18470 19356 18522
rect 19380 18470 19394 18522
rect 19394 18470 19406 18522
rect 19406 18470 19436 18522
rect 19460 18470 19470 18522
rect 19470 18470 19516 18522
rect 19220 18468 19276 18470
rect 19300 18468 19356 18470
rect 19380 18468 19436 18470
rect 19460 18468 19516 18470
rect 19220 17434 19276 17436
rect 19300 17434 19356 17436
rect 19380 17434 19436 17436
rect 19460 17434 19516 17436
rect 19220 17382 19266 17434
rect 19266 17382 19276 17434
rect 19300 17382 19330 17434
rect 19330 17382 19342 17434
rect 19342 17382 19356 17434
rect 19380 17382 19394 17434
rect 19394 17382 19406 17434
rect 19406 17382 19436 17434
rect 19460 17382 19470 17434
rect 19470 17382 19516 17434
rect 19220 17380 19276 17382
rect 19300 17380 19356 17382
rect 19380 17380 19436 17382
rect 19460 17380 19516 17382
rect 16220 10362 16276 10364
rect 16300 10362 16356 10364
rect 16380 10362 16436 10364
rect 16460 10362 16516 10364
rect 16220 10310 16266 10362
rect 16266 10310 16276 10362
rect 16300 10310 16330 10362
rect 16330 10310 16342 10362
rect 16342 10310 16356 10362
rect 16380 10310 16394 10362
rect 16394 10310 16406 10362
rect 16406 10310 16436 10362
rect 16460 10310 16470 10362
rect 16470 10310 16516 10362
rect 16220 10308 16276 10310
rect 16300 10308 16356 10310
rect 16380 10308 16436 10310
rect 16460 10308 16516 10310
rect 13220 4378 13276 4380
rect 13300 4378 13356 4380
rect 13380 4378 13436 4380
rect 13460 4378 13516 4380
rect 13220 4326 13266 4378
rect 13266 4326 13276 4378
rect 13300 4326 13330 4378
rect 13330 4326 13342 4378
rect 13342 4326 13356 4378
rect 13380 4326 13394 4378
rect 13394 4326 13406 4378
rect 13406 4326 13436 4378
rect 13460 4326 13470 4378
rect 13470 4326 13516 4378
rect 13220 4324 13276 4326
rect 13300 4324 13356 4326
rect 13380 4324 13436 4326
rect 13460 4324 13516 4326
rect 13220 3290 13276 3292
rect 13300 3290 13356 3292
rect 13380 3290 13436 3292
rect 13460 3290 13516 3292
rect 13220 3238 13266 3290
rect 13266 3238 13276 3290
rect 13300 3238 13330 3290
rect 13330 3238 13342 3290
rect 13342 3238 13356 3290
rect 13380 3238 13394 3290
rect 13394 3238 13406 3290
rect 13406 3238 13436 3290
rect 13460 3238 13470 3290
rect 13470 3238 13516 3290
rect 13220 3236 13276 3238
rect 13300 3236 13356 3238
rect 13380 3236 13436 3238
rect 13460 3236 13516 3238
rect 16220 9274 16276 9276
rect 16300 9274 16356 9276
rect 16380 9274 16436 9276
rect 16460 9274 16516 9276
rect 16220 9222 16266 9274
rect 16266 9222 16276 9274
rect 16300 9222 16330 9274
rect 16330 9222 16342 9274
rect 16342 9222 16356 9274
rect 16380 9222 16394 9274
rect 16394 9222 16406 9274
rect 16406 9222 16436 9274
rect 16460 9222 16470 9274
rect 16470 9222 16516 9274
rect 16220 9220 16276 9222
rect 16300 9220 16356 9222
rect 16380 9220 16436 9222
rect 16460 9220 16516 9222
rect 19220 16346 19276 16348
rect 19300 16346 19356 16348
rect 19380 16346 19436 16348
rect 19460 16346 19516 16348
rect 19220 16294 19266 16346
rect 19266 16294 19276 16346
rect 19300 16294 19330 16346
rect 19330 16294 19342 16346
rect 19342 16294 19356 16346
rect 19380 16294 19394 16346
rect 19394 16294 19406 16346
rect 19406 16294 19436 16346
rect 19460 16294 19470 16346
rect 19470 16294 19516 16346
rect 19220 16292 19276 16294
rect 19300 16292 19356 16294
rect 19380 16292 19436 16294
rect 19460 16292 19516 16294
rect 19220 15258 19276 15260
rect 19300 15258 19356 15260
rect 19380 15258 19436 15260
rect 19460 15258 19516 15260
rect 19220 15206 19266 15258
rect 19266 15206 19276 15258
rect 19300 15206 19330 15258
rect 19330 15206 19342 15258
rect 19342 15206 19356 15258
rect 19380 15206 19394 15258
rect 19394 15206 19406 15258
rect 19406 15206 19436 15258
rect 19460 15206 19470 15258
rect 19470 15206 19516 15258
rect 19220 15204 19276 15206
rect 19300 15204 19356 15206
rect 19380 15204 19436 15206
rect 19460 15204 19516 15206
rect 20442 21120 20498 21176
rect 19220 14170 19276 14172
rect 19300 14170 19356 14172
rect 19380 14170 19436 14172
rect 19460 14170 19516 14172
rect 19220 14118 19266 14170
rect 19266 14118 19276 14170
rect 19300 14118 19330 14170
rect 19330 14118 19342 14170
rect 19342 14118 19356 14170
rect 19380 14118 19394 14170
rect 19394 14118 19406 14170
rect 19406 14118 19436 14170
rect 19460 14118 19470 14170
rect 19470 14118 19516 14170
rect 19220 14116 19276 14118
rect 19300 14116 19356 14118
rect 19380 14116 19436 14118
rect 19460 14116 19516 14118
rect 19220 13082 19276 13084
rect 19300 13082 19356 13084
rect 19380 13082 19436 13084
rect 19460 13082 19516 13084
rect 19220 13030 19266 13082
rect 19266 13030 19276 13082
rect 19300 13030 19330 13082
rect 19330 13030 19342 13082
rect 19342 13030 19356 13082
rect 19380 13030 19394 13082
rect 19394 13030 19406 13082
rect 19406 13030 19436 13082
rect 19460 13030 19470 13082
rect 19470 13030 19516 13082
rect 19220 13028 19276 13030
rect 19300 13028 19356 13030
rect 19380 13028 19436 13030
rect 19460 13028 19516 13030
rect 19220 11994 19276 11996
rect 19300 11994 19356 11996
rect 19380 11994 19436 11996
rect 19460 11994 19516 11996
rect 19220 11942 19266 11994
rect 19266 11942 19276 11994
rect 19300 11942 19330 11994
rect 19330 11942 19342 11994
rect 19342 11942 19356 11994
rect 19380 11942 19394 11994
rect 19394 11942 19406 11994
rect 19406 11942 19436 11994
rect 19460 11942 19470 11994
rect 19470 11942 19516 11994
rect 19220 11940 19276 11942
rect 19300 11940 19356 11942
rect 19380 11940 19436 11942
rect 19460 11940 19516 11942
rect 19220 10906 19276 10908
rect 19300 10906 19356 10908
rect 19380 10906 19436 10908
rect 19460 10906 19516 10908
rect 19220 10854 19266 10906
rect 19266 10854 19276 10906
rect 19300 10854 19330 10906
rect 19330 10854 19342 10906
rect 19342 10854 19356 10906
rect 19380 10854 19394 10906
rect 19394 10854 19406 10906
rect 19406 10854 19436 10906
rect 19460 10854 19470 10906
rect 19470 10854 19516 10906
rect 19220 10852 19276 10854
rect 19300 10852 19356 10854
rect 19380 10852 19436 10854
rect 19460 10852 19516 10854
rect 19220 9818 19276 9820
rect 19300 9818 19356 9820
rect 19380 9818 19436 9820
rect 19460 9818 19516 9820
rect 19220 9766 19266 9818
rect 19266 9766 19276 9818
rect 19300 9766 19330 9818
rect 19330 9766 19342 9818
rect 19342 9766 19356 9818
rect 19380 9766 19394 9818
rect 19394 9766 19406 9818
rect 19406 9766 19436 9818
rect 19460 9766 19470 9818
rect 19470 9766 19516 9818
rect 19220 9764 19276 9766
rect 19300 9764 19356 9766
rect 19380 9764 19436 9766
rect 19460 9764 19516 9766
rect 16220 8186 16276 8188
rect 16300 8186 16356 8188
rect 16380 8186 16436 8188
rect 16460 8186 16516 8188
rect 16220 8134 16266 8186
rect 16266 8134 16276 8186
rect 16300 8134 16330 8186
rect 16330 8134 16342 8186
rect 16342 8134 16356 8186
rect 16380 8134 16394 8186
rect 16394 8134 16406 8186
rect 16406 8134 16436 8186
rect 16460 8134 16470 8186
rect 16470 8134 16516 8186
rect 16220 8132 16276 8134
rect 16300 8132 16356 8134
rect 16380 8132 16436 8134
rect 16460 8132 16516 8134
rect 16220 7098 16276 7100
rect 16300 7098 16356 7100
rect 16380 7098 16436 7100
rect 16460 7098 16516 7100
rect 16220 7046 16266 7098
rect 16266 7046 16276 7098
rect 16300 7046 16330 7098
rect 16330 7046 16342 7098
rect 16342 7046 16356 7098
rect 16380 7046 16394 7098
rect 16394 7046 16406 7098
rect 16406 7046 16436 7098
rect 16460 7046 16470 7098
rect 16470 7046 16516 7098
rect 16220 7044 16276 7046
rect 16300 7044 16356 7046
rect 16380 7044 16436 7046
rect 16460 7044 16516 7046
rect 16220 6010 16276 6012
rect 16300 6010 16356 6012
rect 16380 6010 16436 6012
rect 16460 6010 16516 6012
rect 16220 5958 16266 6010
rect 16266 5958 16276 6010
rect 16300 5958 16330 6010
rect 16330 5958 16342 6010
rect 16342 5958 16356 6010
rect 16380 5958 16394 6010
rect 16394 5958 16406 6010
rect 16406 5958 16436 6010
rect 16460 5958 16470 6010
rect 16470 5958 16516 6010
rect 16220 5956 16276 5958
rect 16300 5956 16356 5958
rect 16380 5956 16436 5958
rect 16460 5956 16516 5958
rect 19220 8730 19276 8732
rect 19300 8730 19356 8732
rect 19380 8730 19436 8732
rect 19460 8730 19516 8732
rect 19220 8678 19266 8730
rect 19266 8678 19276 8730
rect 19300 8678 19330 8730
rect 19330 8678 19342 8730
rect 19342 8678 19356 8730
rect 19380 8678 19394 8730
rect 19394 8678 19406 8730
rect 19406 8678 19436 8730
rect 19460 8678 19470 8730
rect 19470 8678 19516 8730
rect 19220 8676 19276 8678
rect 19300 8676 19356 8678
rect 19380 8676 19436 8678
rect 19460 8676 19516 8678
rect 20810 10240 20866 10296
rect 19220 7642 19276 7644
rect 19300 7642 19356 7644
rect 19380 7642 19436 7644
rect 19460 7642 19516 7644
rect 19220 7590 19266 7642
rect 19266 7590 19276 7642
rect 19300 7590 19330 7642
rect 19330 7590 19342 7642
rect 19342 7590 19356 7642
rect 19380 7590 19394 7642
rect 19394 7590 19406 7642
rect 19406 7590 19436 7642
rect 19460 7590 19470 7642
rect 19470 7590 19516 7642
rect 19220 7588 19276 7590
rect 19300 7588 19356 7590
rect 19380 7588 19436 7590
rect 19460 7588 19516 7590
rect 19220 6554 19276 6556
rect 19300 6554 19356 6556
rect 19380 6554 19436 6556
rect 19460 6554 19516 6556
rect 19220 6502 19266 6554
rect 19266 6502 19276 6554
rect 19300 6502 19330 6554
rect 19330 6502 19342 6554
rect 19342 6502 19356 6554
rect 19380 6502 19394 6554
rect 19394 6502 19406 6554
rect 19406 6502 19436 6554
rect 19460 6502 19470 6554
rect 19470 6502 19516 6554
rect 19220 6500 19276 6502
rect 19300 6500 19356 6502
rect 19380 6500 19436 6502
rect 19460 6500 19516 6502
rect 19220 5466 19276 5468
rect 19300 5466 19356 5468
rect 19380 5466 19436 5468
rect 19460 5466 19516 5468
rect 19220 5414 19266 5466
rect 19266 5414 19276 5466
rect 19300 5414 19330 5466
rect 19330 5414 19342 5466
rect 19342 5414 19356 5466
rect 19380 5414 19394 5466
rect 19394 5414 19406 5466
rect 19406 5414 19436 5466
rect 19460 5414 19470 5466
rect 19470 5414 19516 5466
rect 19220 5412 19276 5414
rect 19300 5412 19356 5414
rect 19380 5412 19436 5414
rect 19460 5412 19516 5414
rect 16220 4922 16276 4924
rect 16300 4922 16356 4924
rect 16380 4922 16436 4924
rect 16460 4922 16516 4924
rect 16220 4870 16266 4922
rect 16266 4870 16276 4922
rect 16300 4870 16330 4922
rect 16330 4870 16342 4922
rect 16342 4870 16356 4922
rect 16380 4870 16394 4922
rect 16394 4870 16406 4922
rect 16406 4870 16436 4922
rect 16460 4870 16470 4922
rect 16470 4870 16516 4922
rect 16220 4868 16276 4870
rect 16300 4868 16356 4870
rect 16380 4868 16436 4870
rect 16460 4868 16516 4870
rect 20810 4800 20866 4856
rect 19220 4378 19276 4380
rect 19300 4378 19356 4380
rect 19380 4378 19436 4380
rect 19460 4378 19516 4380
rect 19220 4326 19266 4378
rect 19266 4326 19276 4378
rect 19300 4326 19330 4378
rect 19330 4326 19342 4378
rect 19342 4326 19356 4378
rect 19380 4326 19394 4378
rect 19394 4326 19406 4378
rect 19406 4326 19436 4378
rect 19460 4326 19470 4378
rect 19470 4326 19516 4378
rect 19220 4324 19276 4326
rect 19300 4324 19356 4326
rect 19380 4324 19436 4326
rect 19460 4324 19516 4326
rect 16220 3834 16276 3836
rect 16300 3834 16356 3836
rect 16380 3834 16436 3836
rect 16460 3834 16516 3836
rect 16220 3782 16266 3834
rect 16266 3782 16276 3834
rect 16300 3782 16330 3834
rect 16330 3782 16342 3834
rect 16342 3782 16356 3834
rect 16380 3782 16394 3834
rect 16394 3782 16406 3834
rect 16406 3782 16436 3834
rect 16460 3782 16470 3834
rect 16470 3782 16516 3834
rect 16220 3780 16276 3782
rect 16300 3780 16356 3782
rect 16380 3780 16436 3782
rect 16460 3780 16516 3782
rect 19220 3290 19276 3292
rect 19300 3290 19356 3292
rect 19380 3290 19436 3292
rect 19460 3290 19516 3292
rect 19220 3238 19266 3290
rect 19266 3238 19276 3290
rect 19300 3238 19330 3290
rect 19330 3238 19342 3290
rect 19342 3238 19356 3290
rect 19380 3238 19394 3290
rect 19394 3238 19406 3290
rect 19406 3238 19436 3290
rect 19460 3238 19470 3290
rect 19470 3238 19516 3290
rect 19220 3236 19276 3238
rect 19300 3236 19356 3238
rect 19380 3236 19436 3238
rect 19460 3236 19516 3238
rect 16220 2746 16276 2748
rect 16300 2746 16356 2748
rect 16380 2746 16436 2748
rect 16460 2746 16516 2748
rect 16220 2694 16266 2746
rect 16266 2694 16276 2746
rect 16300 2694 16330 2746
rect 16330 2694 16342 2746
rect 16342 2694 16356 2746
rect 16380 2694 16394 2746
rect 16394 2694 16406 2746
rect 16406 2694 16436 2746
rect 16460 2694 16470 2746
rect 16470 2694 16516 2746
rect 16220 2692 16276 2694
rect 16300 2692 16356 2694
rect 16380 2692 16436 2694
rect 16460 2692 16516 2694
rect 13220 2202 13276 2204
rect 13300 2202 13356 2204
rect 13380 2202 13436 2204
rect 13460 2202 13516 2204
rect 13220 2150 13266 2202
rect 13266 2150 13276 2202
rect 13300 2150 13330 2202
rect 13330 2150 13342 2202
rect 13342 2150 13356 2202
rect 13380 2150 13394 2202
rect 13394 2150 13406 2202
rect 13406 2150 13436 2202
rect 13460 2150 13470 2202
rect 13470 2150 13516 2202
rect 13220 2148 13276 2150
rect 13300 2148 13356 2150
rect 13380 2148 13436 2150
rect 13460 2148 13516 2150
rect 19220 2202 19276 2204
rect 19300 2202 19356 2204
rect 19380 2202 19436 2204
rect 19460 2202 19516 2204
rect 19220 2150 19266 2202
rect 19266 2150 19276 2202
rect 19300 2150 19330 2202
rect 19330 2150 19342 2202
rect 19342 2150 19356 2202
rect 19380 2150 19394 2202
rect 19394 2150 19406 2202
rect 19406 2150 19436 2202
rect 19460 2150 19470 2202
rect 19470 2150 19516 2202
rect 19220 2148 19276 2150
rect 19300 2148 19356 2150
rect 19380 2148 19436 2150
rect 19460 2148 19516 2150
<< metal3 >>
rect 0 21858 800 21888
rect 3601 21858 3667 21861
rect 0 21856 3667 21858
rect 0 21800 3606 21856
rect 3662 21800 3667 21856
rect 0 21798 3667 21800
rect 0 21768 800 21798
rect 3601 21795 3667 21798
rect 7210 21792 7526 21793
rect 7210 21728 7216 21792
rect 7280 21728 7296 21792
rect 7360 21728 7376 21792
rect 7440 21728 7456 21792
rect 7520 21728 7526 21792
rect 7210 21727 7526 21728
rect 13210 21792 13526 21793
rect 13210 21728 13216 21792
rect 13280 21728 13296 21792
rect 13360 21728 13376 21792
rect 13440 21728 13456 21792
rect 13520 21728 13526 21792
rect 13210 21727 13526 21728
rect 19210 21792 19526 21793
rect 19210 21728 19216 21792
rect 19280 21728 19296 21792
rect 19360 21728 19376 21792
rect 19440 21728 19456 21792
rect 19520 21728 19526 21792
rect 19210 21727 19526 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 10210 21248 10526 21249
rect 10210 21184 10216 21248
rect 10280 21184 10296 21248
rect 10360 21184 10376 21248
rect 10440 21184 10456 21248
rect 10520 21184 10526 21248
rect 10210 21183 10526 21184
rect 16210 21248 16526 21249
rect 16210 21184 16216 21248
rect 16280 21184 16296 21248
rect 16360 21184 16376 21248
rect 16440 21184 16456 21248
rect 16520 21184 16526 21248
rect 16210 21183 16526 21184
rect 20437 21178 20503 21181
rect 21146 21178 21946 21208
rect 20437 21176 21946 21178
rect 20437 21120 20442 21176
rect 20498 21120 21946 21176
rect 20437 21118 21946 21120
rect 20437 21115 20503 21118
rect 21146 21088 21946 21118
rect 7210 20704 7526 20705
rect 7210 20640 7216 20704
rect 7280 20640 7296 20704
rect 7360 20640 7376 20704
rect 7440 20640 7456 20704
rect 7520 20640 7526 20704
rect 7210 20639 7526 20640
rect 13210 20704 13526 20705
rect 13210 20640 13216 20704
rect 13280 20640 13296 20704
rect 13360 20640 13376 20704
rect 13440 20640 13456 20704
rect 13520 20640 13526 20704
rect 13210 20639 13526 20640
rect 19210 20704 19526 20705
rect 19210 20640 19216 20704
rect 19280 20640 19296 20704
rect 19360 20640 19376 20704
rect 19440 20640 19456 20704
rect 19520 20640 19526 20704
rect 19210 20639 19526 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 10210 20160 10526 20161
rect 10210 20096 10216 20160
rect 10280 20096 10296 20160
rect 10360 20096 10376 20160
rect 10440 20096 10456 20160
rect 10520 20096 10526 20160
rect 10210 20095 10526 20096
rect 16210 20160 16526 20161
rect 16210 20096 16216 20160
rect 16280 20096 16296 20160
rect 16360 20096 16376 20160
rect 16440 20096 16456 20160
rect 16520 20096 16526 20160
rect 16210 20095 16526 20096
rect 7210 19616 7526 19617
rect 7210 19552 7216 19616
rect 7280 19552 7296 19616
rect 7360 19552 7376 19616
rect 7440 19552 7456 19616
rect 7520 19552 7526 19616
rect 7210 19551 7526 19552
rect 13210 19616 13526 19617
rect 13210 19552 13216 19616
rect 13280 19552 13296 19616
rect 13360 19552 13376 19616
rect 13440 19552 13456 19616
rect 13520 19552 13526 19616
rect 13210 19551 13526 19552
rect 19210 19616 19526 19617
rect 19210 19552 19216 19616
rect 19280 19552 19296 19616
rect 19360 19552 19376 19616
rect 19440 19552 19456 19616
rect 19520 19552 19526 19616
rect 19210 19551 19526 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 10210 19072 10526 19073
rect 10210 19008 10216 19072
rect 10280 19008 10296 19072
rect 10360 19008 10376 19072
rect 10440 19008 10456 19072
rect 10520 19008 10526 19072
rect 10210 19007 10526 19008
rect 16210 19072 16526 19073
rect 16210 19008 16216 19072
rect 16280 19008 16296 19072
rect 16360 19008 16376 19072
rect 16440 19008 16456 19072
rect 16520 19008 16526 19072
rect 16210 19007 16526 19008
rect 7210 18528 7526 18529
rect 7210 18464 7216 18528
rect 7280 18464 7296 18528
rect 7360 18464 7376 18528
rect 7440 18464 7456 18528
rect 7520 18464 7526 18528
rect 7210 18463 7526 18464
rect 13210 18528 13526 18529
rect 13210 18464 13216 18528
rect 13280 18464 13296 18528
rect 13360 18464 13376 18528
rect 13440 18464 13456 18528
rect 13520 18464 13526 18528
rect 13210 18463 13526 18464
rect 19210 18528 19526 18529
rect 19210 18464 19216 18528
rect 19280 18464 19296 18528
rect 19360 18464 19376 18528
rect 19440 18464 19456 18528
rect 19520 18464 19526 18528
rect 19210 18463 19526 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 10210 17984 10526 17985
rect 10210 17920 10216 17984
rect 10280 17920 10296 17984
rect 10360 17920 10376 17984
rect 10440 17920 10456 17984
rect 10520 17920 10526 17984
rect 10210 17919 10526 17920
rect 16210 17984 16526 17985
rect 16210 17920 16216 17984
rect 16280 17920 16296 17984
rect 16360 17920 16376 17984
rect 16440 17920 16456 17984
rect 16520 17920 16526 17984
rect 16210 17919 16526 17920
rect 7210 17440 7526 17441
rect 7210 17376 7216 17440
rect 7280 17376 7296 17440
rect 7360 17376 7376 17440
rect 7440 17376 7456 17440
rect 7520 17376 7526 17440
rect 7210 17375 7526 17376
rect 13210 17440 13526 17441
rect 13210 17376 13216 17440
rect 13280 17376 13296 17440
rect 13360 17376 13376 17440
rect 13440 17376 13456 17440
rect 13520 17376 13526 17440
rect 13210 17375 13526 17376
rect 19210 17440 19526 17441
rect 19210 17376 19216 17440
rect 19280 17376 19296 17440
rect 19360 17376 19376 17440
rect 19440 17376 19456 17440
rect 19520 17376 19526 17440
rect 19210 17375 19526 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 10210 16896 10526 16897
rect 10210 16832 10216 16896
rect 10280 16832 10296 16896
rect 10360 16832 10376 16896
rect 10440 16832 10456 16896
rect 10520 16832 10526 16896
rect 10210 16831 10526 16832
rect 16210 16896 16526 16897
rect 16210 16832 16216 16896
rect 16280 16832 16296 16896
rect 16360 16832 16376 16896
rect 16440 16832 16456 16896
rect 16520 16832 16526 16896
rect 16210 16831 16526 16832
rect 0 16418 800 16448
rect 933 16418 999 16421
rect 0 16416 999 16418
rect 0 16360 938 16416
rect 994 16360 999 16416
rect 0 16358 999 16360
rect 0 16328 800 16358
rect 933 16355 999 16358
rect 7210 16352 7526 16353
rect 7210 16288 7216 16352
rect 7280 16288 7296 16352
rect 7360 16288 7376 16352
rect 7440 16288 7456 16352
rect 7520 16288 7526 16352
rect 7210 16287 7526 16288
rect 13210 16352 13526 16353
rect 13210 16288 13216 16352
rect 13280 16288 13296 16352
rect 13360 16288 13376 16352
rect 13440 16288 13456 16352
rect 13520 16288 13526 16352
rect 13210 16287 13526 16288
rect 19210 16352 19526 16353
rect 19210 16288 19216 16352
rect 19280 16288 19296 16352
rect 19360 16288 19376 16352
rect 19440 16288 19456 16352
rect 19520 16288 19526 16352
rect 19210 16287 19526 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 10210 15808 10526 15809
rect 10210 15744 10216 15808
rect 10280 15744 10296 15808
rect 10360 15744 10376 15808
rect 10440 15744 10456 15808
rect 10520 15744 10526 15808
rect 10210 15743 10526 15744
rect 16210 15808 16526 15809
rect 16210 15744 16216 15808
rect 16280 15744 16296 15808
rect 16360 15744 16376 15808
rect 16440 15744 16456 15808
rect 16520 15744 16526 15808
rect 16210 15743 16526 15744
rect 17033 15738 17099 15741
rect 21146 15738 21946 15768
rect 17033 15736 21946 15738
rect 17033 15680 17038 15736
rect 17094 15680 21946 15736
rect 17033 15678 21946 15680
rect 17033 15675 17099 15678
rect 21146 15648 21946 15678
rect 7210 15264 7526 15265
rect 7210 15200 7216 15264
rect 7280 15200 7296 15264
rect 7360 15200 7376 15264
rect 7440 15200 7456 15264
rect 7520 15200 7526 15264
rect 7210 15199 7526 15200
rect 13210 15264 13526 15265
rect 13210 15200 13216 15264
rect 13280 15200 13296 15264
rect 13360 15200 13376 15264
rect 13440 15200 13456 15264
rect 13520 15200 13526 15264
rect 13210 15199 13526 15200
rect 19210 15264 19526 15265
rect 19210 15200 19216 15264
rect 19280 15200 19296 15264
rect 19360 15200 19376 15264
rect 19440 15200 19456 15264
rect 19520 15200 19526 15264
rect 19210 15199 19526 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 10210 14720 10526 14721
rect 10210 14656 10216 14720
rect 10280 14656 10296 14720
rect 10360 14656 10376 14720
rect 10440 14656 10456 14720
rect 10520 14656 10526 14720
rect 10210 14655 10526 14656
rect 16210 14720 16526 14721
rect 16210 14656 16216 14720
rect 16280 14656 16296 14720
rect 16360 14656 16376 14720
rect 16440 14656 16456 14720
rect 16520 14656 16526 14720
rect 16210 14655 16526 14656
rect 7210 14176 7526 14177
rect 7210 14112 7216 14176
rect 7280 14112 7296 14176
rect 7360 14112 7376 14176
rect 7440 14112 7456 14176
rect 7520 14112 7526 14176
rect 7210 14111 7526 14112
rect 13210 14176 13526 14177
rect 13210 14112 13216 14176
rect 13280 14112 13296 14176
rect 13360 14112 13376 14176
rect 13440 14112 13456 14176
rect 13520 14112 13526 14176
rect 13210 14111 13526 14112
rect 19210 14176 19526 14177
rect 19210 14112 19216 14176
rect 19280 14112 19296 14176
rect 19360 14112 19376 14176
rect 19440 14112 19456 14176
rect 19520 14112 19526 14176
rect 19210 14111 19526 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 10210 13632 10526 13633
rect 10210 13568 10216 13632
rect 10280 13568 10296 13632
rect 10360 13568 10376 13632
rect 10440 13568 10456 13632
rect 10520 13568 10526 13632
rect 10210 13567 10526 13568
rect 16210 13632 16526 13633
rect 16210 13568 16216 13632
rect 16280 13568 16296 13632
rect 16360 13568 16376 13632
rect 16440 13568 16456 13632
rect 16520 13568 16526 13632
rect 16210 13567 16526 13568
rect 7210 13088 7526 13089
rect 7210 13024 7216 13088
rect 7280 13024 7296 13088
rect 7360 13024 7376 13088
rect 7440 13024 7456 13088
rect 7520 13024 7526 13088
rect 7210 13023 7526 13024
rect 13210 13088 13526 13089
rect 13210 13024 13216 13088
rect 13280 13024 13296 13088
rect 13360 13024 13376 13088
rect 13440 13024 13456 13088
rect 13520 13024 13526 13088
rect 13210 13023 13526 13024
rect 19210 13088 19526 13089
rect 19210 13024 19216 13088
rect 19280 13024 19296 13088
rect 19360 13024 19376 13088
rect 19440 13024 19456 13088
rect 19520 13024 19526 13088
rect 19210 13023 19526 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 10210 12544 10526 12545
rect 10210 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10526 12544
rect 10210 12479 10526 12480
rect 16210 12544 16526 12545
rect 16210 12480 16216 12544
rect 16280 12480 16296 12544
rect 16360 12480 16376 12544
rect 16440 12480 16456 12544
rect 16520 12480 16526 12544
rect 16210 12479 16526 12480
rect 7210 12000 7526 12001
rect 7210 11936 7216 12000
rect 7280 11936 7296 12000
rect 7360 11936 7376 12000
rect 7440 11936 7456 12000
rect 7520 11936 7526 12000
rect 7210 11935 7526 11936
rect 13210 12000 13526 12001
rect 13210 11936 13216 12000
rect 13280 11936 13296 12000
rect 13360 11936 13376 12000
rect 13440 11936 13456 12000
rect 13520 11936 13526 12000
rect 13210 11935 13526 11936
rect 19210 12000 19526 12001
rect 19210 11936 19216 12000
rect 19280 11936 19296 12000
rect 19360 11936 19376 12000
rect 19440 11936 19456 12000
rect 19520 11936 19526 12000
rect 19210 11935 19526 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 10210 11456 10526 11457
rect 10210 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10526 11456
rect 10210 11391 10526 11392
rect 16210 11456 16526 11457
rect 16210 11392 16216 11456
rect 16280 11392 16296 11456
rect 16360 11392 16376 11456
rect 16440 11392 16456 11456
rect 16520 11392 16526 11456
rect 16210 11391 16526 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 7210 10912 7526 10913
rect 7210 10848 7216 10912
rect 7280 10848 7296 10912
rect 7360 10848 7376 10912
rect 7440 10848 7456 10912
rect 7520 10848 7526 10912
rect 7210 10847 7526 10848
rect 13210 10912 13526 10913
rect 13210 10848 13216 10912
rect 13280 10848 13296 10912
rect 13360 10848 13376 10912
rect 13440 10848 13456 10912
rect 13520 10848 13526 10912
rect 13210 10847 13526 10848
rect 19210 10912 19526 10913
rect 19210 10848 19216 10912
rect 19280 10848 19296 10912
rect 19360 10848 19376 10912
rect 19440 10848 19456 10912
rect 19520 10848 19526 10912
rect 19210 10847 19526 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 10210 10368 10526 10369
rect 10210 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10526 10368
rect 10210 10303 10526 10304
rect 16210 10368 16526 10369
rect 16210 10304 16216 10368
rect 16280 10304 16296 10368
rect 16360 10304 16376 10368
rect 16440 10304 16456 10368
rect 16520 10304 16526 10368
rect 16210 10303 16526 10304
rect 20805 10298 20871 10301
rect 21146 10298 21946 10328
rect 20805 10296 21946 10298
rect 20805 10240 20810 10296
rect 20866 10240 21946 10296
rect 20805 10238 21946 10240
rect 20805 10235 20871 10238
rect 21146 10208 21946 10238
rect 7210 9824 7526 9825
rect 7210 9760 7216 9824
rect 7280 9760 7296 9824
rect 7360 9760 7376 9824
rect 7440 9760 7456 9824
rect 7520 9760 7526 9824
rect 7210 9759 7526 9760
rect 13210 9824 13526 9825
rect 13210 9760 13216 9824
rect 13280 9760 13296 9824
rect 13360 9760 13376 9824
rect 13440 9760 13456 9824
rect 13520 9760 13526 9824
rect 13210 9759 13526 9760
rect 19210 9824 19526 9825
rect 19210 9760 19216 9824
rect 19280 9760 19296 9824
rect 19360 9760 19376 9824
rect 19440 9760 19456 9824
rect 19520 9760 19526 9824
rect 19210 9759 19526 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 10210 9280 10526 9281
rect 10210 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10526 9280
rect 10210 9215 10526 9216
rect 16210 9280 16526 9281
rect 16210 9216 16216 9280
rect 16280 9216 16296 9280
rect 16360 9216 16376 9280
rect 16440 9216 16456 9280
rect 16520 9216 16526 9280
rect 16210 9215 16526 9216
rect 7210 8736 7526 8737
rect 7210 8672 7216 8736
rect 7280 8672 7296 8736
rect 7360 8672 7376 8736
rect 7440 8672 7456 8736
rect 7520 8672 7526 8736
rect 7210 8671 7526 8672
rect 13210 8736 13526 8737
rect 13210 8672 13216 8736
rect 13280 8672 13296 8736
rect 13360 8672 13376 8736
rect 13440 8672 13456 8736
rect 13520 8672 13526 8736
rect 13210 8671 13526 8672
rect 19210 8736 19526 8737
rect 19210 8672 19216 8736
rect 19280 8672 19296 8736
rect 19360 8672 19376 8736
rect 19440 8672 19456 8736
rect 19520 8672 19526 8736
rect 19210 8671 19526 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 10210 8192 10526 8193
rect 10210 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10526 8192
rect 10210 8127 10526 8128
rect 16210 8192 16526 8193
rect 16210 8128 16216 8192
rect 16280 8128 16296 8192
rect 16360 8128 16376 8192
rect 16440 8128 16456 8192
rect 16520 8128 16526 8192
rect 16210 8127 16526 8128
rect 7210 7648 7526 7649
rect 7210 7584 7216 7648
rect 7280 7584 7296 7648
rect 7360 7584 7376 7648
rect 7440 7584 7456 7648
rect 7520 7584 7526 7648
rect 7210 7583 7526 7584
rect 13210 7648 13526 7649
rect 13210 7584 13216 7648
rect 13280 7584 13296 7648
rect 13360 7584 13376 7648
rect 13440 7584 13456 7648
rect 13520 7584 13526 7648
rect 13210 7583 13526 7584
rect 19210 7648 19526 7649
rect 19210 7584 19216 7648
rect 19280 7584 19296 7648
rect 19360 7584 19376 7648
rect 19440 7584 19456 7648
rect 19520 7584 19526 7648
rect 19210 7583 19526 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 10210 7104 10526 7105
rect 10210 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10526 7104
rect 10210 7039 10526 7040
rect 16210 7104 16526 7105
rect 16210 7040 16216 7104
rect 16280 7040 16296 7104
rect 16360 7040 16376 7104
rect 16440 7040 16456 7104
rect 16520 7040 16526 7104
rect 16210 7039 16526 7040
rect 7210 6560 7526 6561
rect 7210 6496 7216 6560
rect 7280 6496 7296 6560
rect 7360 6496 7376 6560
rect 7440 6496 7456 6560
rect 7520 6496 7526 6560
rect 7210 6495 7526 6496
rect 13210 6560 13526 6561
rect 13210 6496 13216 6560
rect 13280 6496 13296 6560
rect 13360 6496 13376 6560
rect 13440 6496 13456 6560
rect 13520 6496 13526 6560
rect 13210 6495 13526 6496
rect 19210 6560 19526 6561
rect 19210 6496 19216 6560
rect 19280 6496 19296 6560
rect 19360 6496 19376 6560
rect 19440 6496 19456 6560
rect 19520 6496 19526 6560
rect 19210 6495 19526 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 10210 6016 10526 6017
rect 10210 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10526 6016
rect 10210 5951 10526 5952
rect 16210 6016 16526 6017
rect 16210 5952 16216 6016
rect 16280 5952 16296 6016
rect 16360 5952 16376 6016
rect 16440 5952 16456 6016
rect 16520 5952 16526 6016
rect 16210 5951 16526 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 7210 5472 7526 5473
rect 7210 5408 7216 5472
rect 7280 5408 7296 5472
rect 7360 5408 7376 5472
rect 7440 5408 7456 5472
rect 7520 5408 7526 5472
rect 7210 5407 7526 5408
rect 13210 5472 13526 5473
rect 13210 5408 13216 5472
rect 13280 5408 13296 5472
rect 13360 5408 13376 5472
rect 13440 5408 13456 5472
rect 13520 5408 13526 5472
rect 13210 5407 13526 5408
rect 19210 5472 19526 5473
rect 19210 5408 19216 5472
rect 19280 5408 19296 5472
rect 19360 5408 19376 5472
rect 19440 5408 19456 5472
rect 19520 5408 19526 5472
rect 19210 5407 19526 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 10210 4928 10526 4929
rect 10210 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10526 4928
rect 10210 4863 10526 4864
rect 16210 4928 16526 4929
rect 16210 4864 16216 4928
rect 16280 4864 16296 4928
rect 16360 4864 16376 4928
rect 16440 4864 16456 4928
rect 16520 4864 16526 4928
rect 16210 4863 16526 4864
rect 20805 4858 20871 4861
rect 21146 4858 21946 4888
rect 20805 4856 21946 4858
rect 20805 4800 20810 4856
rect 20866 4800 21946 4856
rect 20805 4798 21946 4800
rect 20805 4795 20871 4798
rect 21146 4768 21946 4798
rect 7210 4384 7526 4385
rect 7210 4320 7216 4384
rect 7280 4320 7296 4384
rect 7360 4320 7376 4384
rect 7440 4320 7456 4384
rect 7520 4320 7526 4384
rect 7210 4319 7526 4320
rect 13210 4384 13526 4385
rect 13210 4320 13216 4384
rect 13280 4320 13296 4384
rect 13360 4320 13376 4384
rect 13440 4320 13456 4384
rect 13520 4320 13526 4384
rect 13210 4319 13526 4320
rect 19210 4384 19526 4385
rect 19210 4320 19216 4384
rect 19280 4320 19296 4384
rect 19360 4320 19376 4384
rect 19440 4320 19456 4384
rect 19520 4320 19526 4384
rect 19210 4319 19526 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 10210 3840 10526 3841
rect 10210 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10526 3840
rect 10210 3775 10526 3776
rect 16210 3840 16526 3841
rect 16210 3776 16216 3840
rect 16280 3776 16296 3840
rect 16360 3776 16376 3840
rect 16440 3776 16456 3840
rect 16520 3776 16526 3840
rect 16210 3775 16526 3776
rect 7210 3296 7526 3297
rect 7210 3232 7216 3296
rect 7280 3232 7296 3296
rect 7360 3232 7376 3296
rect 7440 3232 7456 3296
rect 7520 3232 7526 3296
rect 7210 3231 7526 3232
rect 13210 3296 13526 3297
rect 13210 3232 13216 3296
rect 13280 3232 13296 3296
rect 13360 3232 13376 3296
rect 13440 3232 13456 3296
rect 13520 3232 13526 3296
rect 13210 3231 13526 3232
rect 19210 3296 19526 3297
rect 19210 3232 19216 3296
rect 19280 3232 19296 3296
rect 19360 3232 19376 3296
rect 19440 3232 19456 3296
rect 19520 3232 19526 3296
rect 19210 3231 19526 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 10210 2752 10526 2753
rect 10210 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10526 2752
rect 10210 2687 10526 2688
rect 16210 2752 16526 2753
rect 16210 2688 16216 2752
rect 16280 2688 16296 2752
rect 16360 2688 16376 2752
rect 16440 2688 16456 2752
rect 16520 2688 16526 2752
rect 16210 2687 16526 2688
rect 7210 2208 7526 2209
rect 7210 2144 7216 2208
rect 7280 2144 7296 2208
rect 7360 2144 7376 2208
rect 7440 2144 7456 2208
rect 7520 2144 7526 2208
rect 7210 2143 7526 2144
rect 13210 2208 13526 2209
rect 13210 2144 13216 2208
rect 13280 2144 13296 2208
rect 13360 2144 13376 2208
rect 13440 2144 13456 2208
rect 13520 2144 13526 2208
rect 13210 2143 13526 2144
rect 19210 2208 19526 2209
rect 19210 2144 19216 2208
rect 19280 2144 19296 2208
rect 19360 2144 19376 2208
rect 19440 2144 19456 2208
rect 19520 2144 19526 2208
rect 19210 2143 19526 2144
<< via3 >>
rect 7216 21788 7280 21792
rect 7216 21732 7220 21788
rect 7220 21732 7276 21788
rect 7276 21732 7280 21788
rect 7216 21728 7280 21732
rect 7296 21788 7360 21792
rect 7296 21732 7300 21788
rect 7300 21732 7356 21788
rect 7356 21732 7360 21788
rect 7296 21728 7360 21732
rect 7376 21788 7440 21792
rect 7376 21732 7380 21788
rect 7380 21732 7436 21788
rect 7436 21732 7440 21788
rect 7376 21728 7440 21732
rect 7456 21788 7520 21792
rect 7456 21732 7460 21788
rect 7460 21732 7516 21788
rect 7516 21732 7520 21788
rect 7456 21728 7520 21732
rect 13216 21788 13280 21792
rect 13216 21732 13220 21788
rect 13220 21732 13276 21788
rect 13276 21732 13280 21788
rect 13216 21728 13280 21732
rect 13296 21788 13360 21792
rect 13296 21732 13300 21788
rect 13300 21732 13356 21788
rect 13356 21732 13360 21788
rect 13296 21728 13360 21732
rect 13376 21788 13440 21792
rect 13376 21732 13380 21788
rect 13380 21732 13436 21788
rect 13436 21732 13440 21788
rect 13376 21728 13440 21732
rect 13456 21788 13520 21792
rect 13456 21732 13460 21788
rect 13460 21732 13516 21788
rect 13516 21732 13520 21788
rect 13456 21728 13520 21732
rect 19216 21788 19280 21792
rect 19216 21732 19220 21788
rect 19220 21732 19276 21788
rect 19276 21732 19280 21788
rect 19216 21728 19280 21732
rect 19296 21788 19360 21792
rect 19296 21732 19300 21788
rect 19300 21732 19356 21788
rect 19356 21732 19360 21788
rect 19296 21728 19360 21732
rect 19376 21788 19440 21792
rect 19376 21732 19380 21788
rect 19380 21732 19436 21788
rect 19436 21732 19440 21788
rect 19376 21728 19440 21732
rect 19456 21788 19520 21792
rect 19456 21732 19460 21788
rect 19460 21732 19516 21788
rect 19516 21732 19520 21788
rect 19456 21728 19520 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 10216 21244 10280 21248
rect 10216 21188 10220 21244
rect 10220 21188 10276 21244
rect 10276 21188 10280 21244
rect 10216 21184 10280 21188
rect 10296 21244 10360 21248
rect 10296 21188 10300 21244
rect 10300 21188 10356 21244
rect 10356 21188 10360 21244
rect 10296 21184 10360 21188
rect 10376 21244 10440 21248
rect 10376 21188 10380 21244
rect 10380 21188 10436 21244
rect 10436 21188 10440 21244
rect 10376 21184 10440 21188
rect 10456 21244 10520 21248
rect 10456 21188 10460 21244
rect 10460 21188 10516 21244
rect 10516 21188 10520 21244
rect 10456 21184 10520 21188
rect 16216 21244 16280 21248
rect 16216 21188 16220 21244
rect 16220 21188 16276 21244
rect 16276 21188 16280 21244
rect 16216 21184 16280 21188
rect 16296 21244 16360 21248
rect 16296 21188 16300 21244
rect 16300 21188 16356 21244
rect 16356 21188 16360 21244
rect 16296 21184 16360 21188
rect 16376 21244 16440 21248
rect 16376 21188 16380 21244
rect 16380 21188 16436 21244
rect 16436 21188 16440 21244
rect 16376 21184 16440 21188
rect 16456 21244 16520 21248
rect 16456 21188 16460 21244
rect 16460 21188 16516 21244
rect 16516 21188 16520 21244
rect 16456 21184 16520 21188
rect 7216 20700 7280 20704
rect 7216 20644 7220 20700
rect 7220 20644 7276 20700
rect 7276 20644 7280 20700
rect 7216 20640 7280 20644
rect 7296 20700 7360 20704
rect 7296 20644 7300 20700
rect 7300 20644 7356 20700
rect 7356 20644 7360 20700
rect 7296 20640 7360 20644
rect 7376 20700 7440 20704
rect 7376 20644 7380 20700
rect 7380 20644 7436 20700
rect 7436 20644 7440 20700
rect 7376 20640 7440 20644
rect 7456 20700 7520 20704
rect 7456 20644 7460 20700
rect 7460 20644 7516 20700
rect 7516 20644 7520 20700
rect 7456 20640 7520 20644
rect 13216 20700 13280 20704
rect 13216 20644 13220 20700
rect 13220 20644 13276 20700
rect 13276 20644 13280 20700
rect 13216 20640 13280 20644
rect 13296 20700 13360 20704
rect 13296 20644 13300 20700
rect 13300 20644 13356 20700
rect 13356 20644 13360 20700
rect 13296 20640 13360 20644
rect 13376 20700 13440 20704
rect 13376 20644 13380 20700
rect 13380 20644 13436 20700
rect 13436 20644 13440 20700
rect 13376 20640 13440 20644
rect 13456 20700 13520 20704
rect 13456 20644 13460 20700
rect 13460 20644 13516 20700
rect 13516 20644 13520 20700
rect 13456 20640 13520 20644
rect 19216 20700 19280 20704
rect 19216 20644 19220 20700
rect 19220 20644 19276 20700
rect 19276 20644 19280 20700
rect 19216 20640 19280 20644
rect 19296 20700 19360 20704
rect 19296 20644 19300 20700
rect 19300 20644 19356 20700
rect 19356 20644 19360 20700
rect 19296 20640 19360 20644
rect 19376 20700 19440 20704
rect 19376 20644 19380 20700
rect 19380 20644 19436 20700
rect 19436 20644 19440 20700
rect 19376 20640 19440 20644
rect 19456 20700 19520 20704
rect 19456 20644 19460 20700
rect 19460 20644 19516 20700
rect 19516 20644 19520 20700
rect 19456 20640 19520 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 10216 20156 10280 20160
rect 10216 20100 10220 20156
rect 10220 20100 10276 20156
rect 10276 20100 10280 20156
rect 10216 20096 10280 20100
rect 10296 20156 10360 20160
rect 10296 20100 10300 20156
rect 10300 20100 10356 20156
rect 10356 20100 10360 20156
rect 10296 20096 10360 20100
rect 10376 20156 10440 20160
rect 10376 20100 10380 20156
rect 10380 20100 10436 20156
rect 10436 20100 10440 20156
rect 10376 20096 10440 20100
rect 10456 20156 10520 20160
rect 10456 20100 10460 20156
rect 10460 20100 10516 20156
rect 10516 20100 10520 20156
rect 10456 20096 10520 20100
rect 16216 20156 16280 20160
rect 16216 20100 16220 20156
rect 16220 20100 16276 20156
rect 16276 20100 16280 20156
rect 16216 20096 16280 20100
rect 16296 20156 16360 20160
rect 16296 20100 16300 20156
rect 16300 20100 16356 20156
rect 16356 20100 16360 20156
rect 16296 20096 16360 20100
rect 16376 20156 16440 20160
rect 16376 20100 16380 20156
rect 16380 20100 16436 20156
rect 16436 20100 16440 20156
rect 16376 20096 16440 20100
rect 16456 20156 16520 20160
rect 16456 20100 16460 20156
rect 16460 20100 16516 20156
rect 16516 20100 16520 20156
rect 16456 20096 16520 20100
rect 7216 19612 7280 19616
rect 7216 19556 7220 19612
rect 7220 19556 7276 19612
rect 7276 19556 7280 19612
rect 7216 19552 7280 19556
rect 7296 19612 7360 19616
rect 7296 19556 7300 19612
rect 7300 19556 7356 19612
rect 7356 19556 7360 19612
rect 7296 19552 7360 19556
rect 7376 19612 7440 19616
rect 7376 19556 7380 19612
rect 7380 19556 7436 19612
rect 7436 19556 7440 19612
rect 7376 19552 7440 19556
rect 7456 19612 7520 19616
rect 7456 19556 7460 19612
rect 7460 19556 7516 19612
rect 7516 19556 7520 19612
rect 7456 19552 7520 19556
rect 13216 19612 13280 19616
rect 13216 19556 13220 19612
rect 13220 19556 13276 19612
rect 13276 19556 13280 19612
rect 13216 19552 13280 19556
rect 13296 19612 13360 19616
rect 13296 19556 13300 19612
rect 13300 19556 13356 19612
rect 13356 19556 13360 19612
rect 13296 19552 13360 19556
rect 13376 19612 13440 19616
rect 13376 19556 13380 19612
rect 13380 19556 13436 19612
rect 13436 19556 13440 19612
rect 13376 19552 13440 19556
rect 13456 19612 13520 19616
rect 13456 19556 13460 19612
rect 13460 19556 13516 19612
rect 13516 19556 13520 19612
rect 13456 19552 13520 19556
rect 19216 19612 19280 19616
rect 19216 19556 19220 19612
rect 19220 19556 19276 19612
rect 19276 19556 19280 19612
rect 19216 19552 19280 19556
rect 19296 19612 19360 19616
rect 19296 19556 19300 19612
rect 19300 19556 19356 19612
rect 19356 19556 19360 19612
rect 19296 19552 19360 19556
rect 19376 19612 19440 19616
rect 19376 19556 19380 19612
rect 19380 19556 19436 19612
rect 19436 19556 19440 19612
rect 19376 19552 19440 19556
rect 19456 19612 19520 19616
rect 19456 19556 19460 19612
rect 19460 19556 19516 19612
rect 19516 19556 19520 19612
rect 19456 19552 19520 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 10216 19068 10280 19072
rect 10216 19012 10220 19068
rect 10220 19012 10276 19068
rect 10276 19012 10280 19068
rect 10216 19008 10280 19012
rect 10296 19068 10360 19072
rect 10296 19012 10300 19068
rect 10300 19012 10356 19068
rect 10356 19012 10360 19068
rect 10296 19008 10360 19012
rect 10376 19068 10440 19072
rect 10376 19012 10380 19068
rect 10380 19012 10436 19068
rect 10436 19012 10440 19068
rect 10376 19008 10440 19012
rect 10456 19068 10520 19072
rect 10456 19012 10460 19068
rect 10460 19012 10516 19068
rect 10516 19012 10520 19068
rect 10456 19008 10520 19012
rect 16216 19068 16280 19072
rect 16216 19012 16220 19068
rect 16220 19012 16276 19068
rect 16276 19012 16280 19068
rect 16216 19008 16280 19012
rect 16296 19068 16360 19072
rect 16296 19012 16300 19068
rect 16300 19012 16356 19068
rect 16356 19012 16360 19068
rect 16296 19008 16360 19012
rect 16376 19068 16440 19072
rect 16376 19012 16380 19068
rect 16380 19012 16436 19068
rect 16436 19012 16440 19068
rect 16376 19008 16440 19012
rect 16456 19068 16520 19072
rect 16456 19012 16460 19068
rect 16460 19012 16516 19068
rect 16516 19012 16520 19068
rect 16456 19008 16520 19012
rect 7216 18524 7280 18528
rect 7216 18468 7220 18524
rect 7220 18468 7276 18524
rect 7276 18468 7280 18524
rect 7216 18464 7280 18468
rect 7296 18524 7360 18528
rect 7296 18468 7300 18524
rect 7300 18468 7356 18524
rect 7356 18468 7360 18524
rect 7296 18464 7360 18468
rect 7376 18524 7440 18528
rect 7376 18468 7380 18524
rect 7380 18468 7436 18524
rect 7436 18468 7440 18524
rect 7376 18464 7440 18468
rect 7456 18524 7520 18528
rect 7456 18468 7460 18524
rect 7460 18468 7516 18524
rect 7516 18468 7520 18524
rect 7456 18464 7520 18468
rect 13216 18524 13280 18528
rect 13216 18468 13220 18524
rect 13220 18468 13276 18524
rect 13276 18468 13280 18524
rect 13216 18464 13280 18468
rect 13296 18524 13360 18528
rect 13296 18468 13300 18524
rect 13300 18468 13356 18524
rect 13356 18468 13360 18524
rect 13296 18464 13360 18468
rect 13376 18524 13440 18528
rect 13376 18468 13380 18524
rect 13380 18468 13436 18524
rect 13436 18468 13440 18524
rect 13376 18464 13440 18468
rect 13456 18524 13520 18528
rect 13456 18468 13460 18524
rect 13460 18468 13516 18524
rect 13516 18468 13520 18524
rect 13456 18464 13520 18468
rect 19216 18524 19280 18528
rect 19216 18468 19220 18524
rect 19220 18468 19276 18524
rect 19276 18468 19280 18524
rect 19216 18464 19280 18468
rect 19296 18524 19360 18528
rect 19296 18468 19300 18524
rect 19300 18468 19356 18524
rect 19356 18468 19360 18524
rect 19296 18464 19360 18468
rect 19376 18524 19440 18528
rect 19376 18468 19380 18524
rect 19380 18468 19436 18524
rect 19436 18468 19440 18524
rect 19376 18464 19440 18468
rect 19456 18524 19520 18528
rect 19456 18468 19460 18524
rect 19460 18468 19516 18524
rect 19516 18468 19520 18524
rect 19456 18464 19520 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 10216 17980 10280 17984
rect 10216 17924 10220 17980
rect 10220 17924 10276 17980
rect 10276 17924 10280 17980
rect 10216 17920 10280 17924
rect 10296 17980 10360 17984
rect 10296 17924 10300 17980
rect 10300 17924 10356 17980
rect 10356 17924 10360 17980
rect 10296 17920 10360 17924
rect 10376 17980 10440 17984
rect 10376 17924 10380 17980
rect 10380 17924 10436 17980
rect 10436 17924 10440 17980
rect 10376 17920 10440 17924
rect 10456 17980 10520 17984
rect 10456 17924 10460 17980
rect 10460 17924 10516 17980
rect 10516 17924 10520 17980
rect 10456 17920 10520 17924
rect 16216 17980 16280 17984
rect 16216 17924 16220 17980
rect 16220 17924 16276 17980
rect 16276 17924 16280 17980
rect 16216 17920 16280 17924
rect 16296 17980 16360 17984
rect 16296 17924 16300 17980
rect 16300 17924 16356 17980
rect 16356 17924 16360 17980
rect 16296 17920 16360 17924
rect 16376 17980 16440 17984
rect 16376 17924 16380 17980
rect 16380 17924 16436 17980
rect 16436 17924 16440 17980
rect 16376 17920 16440 17924
rect 16456 17980 16520 17984
rect 16456 17924 16460 17980
rect 16460 17924 16516 17980
rect 16516 17924 16520 17980
rect 16456 17920 16520 17924
rect 7216 17436 7280 17440
rect 7216 17380 7220 17436
rect 7220 17380 7276 17436
rect 7276 17380 7280 17436
rect 7216 17376 7280 17380
rect 7296 17436 7360 17440
rect 7296 17380 7300 17436
rect 7300 17380 7356 17436
rect 7356 17380 7360 17436
rect 7296 17376 7360 17380
rect 7376 17436 7440 17440
rect 7376 17380 7380 17436
rect 7380 17380 7436 17436
rect 7436 17380 7440 17436
rect 7376 17376 7440 17380
rect 7456 17436 7520 17440
rect 7456 17380 7460 17436
rect 7460 17380 7516 17436
rect 7516 17380 7520 17436
rect 7456 17376 7520 17380
rect 13216 17436 13280 17440
rect 13216 17380 13220 17436
rect 13220 17380 13276 17436
rect 13276 17380 13280 17436
rect 13216 17376 13280 17380
rect 13296 17436 13360 17440
rect 13296 17380 13300 17436
rect 13300 17380 13356 17436
rect 13356 17380 13360 17436
rect 13296 17376 13360 17380
rect 13376 17436 13440 17440
rect 13376 17380 13380 17436
rect 13380 17380 13436 17436
rect 13436 17380 13440 17436
rect 13376 17376 13440 17380
rect 13456 17436 13520 17440
rect 13456 17380 13460 17436
rect 13460 17380 13516 17436
rect 13516 17380 13520 17436
rect 13456 17376 13520 17380
rect 19216 17436 19280 17440
rect 19216 17380 19220 17436
rect 19220 17380 19276 17436
rect 19276 17380 19280 17436
rect 19216 17376 19280 17380
rect 19296 17436 19360 17440
rect 19296 17380 19300 17436
rect 19300 17380 19356 17436
rect 19356 17380 19360 17436
rect 19296 17376 19360 17380
rect 19376 17436 19440 17440
rect 19376 17380 19380 17436
rect 19380 17380 19436 17436
rect 19436 17380 19440 17436
rect 19376 17376 19440 17380
rect 19456 17436 19520 17440
rect 19456 17380 19460 17436
rect 19460 17380 19516 17436
rect 19516 17380 19520 17436
rect 19456 17376 19520 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 10216 16892 10280 16896
rect 10216 16836 10220 16892
rect 10220 16836 10276 16892
rect 10276 16836 10280 16892
rect 10216 16832 10280 16836
rect 10296 16892 10360 16896
rect 10296 16836 10300 16892
rect 10300 16836 10356 16892
rect 10356 16836 10360 16892
rect 10296 16832 10360 16836
rect 10376 16892 10440 16896
rect 10376 16836 10380 16892
rect 10380 16836 10436 16892
rect 10436 16836 10440 16892
rect 10376 16832 10440 16836
rect 10456 16892 10520 16896
rect 10456 16836 10460 16892
rect 10460 16836 10516 16892
rect 10516 16836 10520 16892
rect 10456 16832 10520 16836
rect 16216 16892 16280 16896
rect 16216 16836 16220 16892
rect 16220 16836 16276 16892
rect 16276 16836 16280 16892
rect 16216 16832 16280 16836
rect 16296 16892 16360 16896
rect 16296 16836 16300 16892
rect 16300 16836 16356 16892
rect 16356 16836 16360 16892
rect 16296 16832 16360 16836
rect 16376 16892 16440 16896
rect 16376 16836 16380 16892
rect 16380 16836 16436 16892
rect 16436 16836 16440 16892
rect 16376 16832 16440 16836
rect 16456 16892 16520 16896
rect 16456 16836 16460 16892
rect 16460 16836 16516 16892
rect 16516 16836 16520 16892
rect 16456 16832 16520 16836
rect 7216 16348 7280 16352
rect 7216 16292 7220 16348
rect 7220 16292 7276 16348
rect 7276 16292 7280 16348
rect 7216 16288 7280 16292
rect 7296 16348 7360 16352
rect 7296 16292 7300 16348
rect 7300 16292 7356 16348
rect 7356 16292 7360 16348
rect 7296 16288 7360 16292
rect 7376 16348 7440 16352
rect 7376 16292 7380 16348
rect 7380 16292 7436 16348
rect 7436 16292 7440 16348
rect 7376 16288 7440 16292
rect 7456 16348 7520 16352
rect 7456 16292 7460 16348
rect 7460 16292 7516 16348
rect 7516 16292 7520 16348
rect 7456 16288 7520 16292
rect 13216 16348 13280 16352
rect 13216 16292 13220 16348
rect 13220 16292 13276 16348
rect 13276 16292 13280 16348
rect 13216 16288 13280 16292
rect 13296 16348 13360 16352
rect 13296 16292 13300 16348
rect 13300 16292 13356 16348
rect 13356 16292 13360 16348
rect 13296 16288 13360 16292
rect 13376 16348 13440 16352
rect 13376 16292 13380 16348
rect 13380 16292 13436 16348
rect 13436 16292 13440 16348
rect 13376 16288 13440 16292
rect 13456 16348 13520 16352
rect 13456 16292 13460 16348
rect 13460 16292 13516 16348
rect 13516 16292 13520 16348
rect 13456 16288 13520 16292
rect 19216 16348 19280 16352
rect 19216 16292 19220 16348
rect 19220 16292 19276 16348
rect 19276 16292 19280 16348
rect 19216 16288 19280 16292
rect 19296 16348 19360 16352
rect 19296 16292 19300 16348
rect 19300 16292 19356 16348
rect 19356 16292 19360 16348
rect 19296 16288 19360 16292
rect 19376 16348 19440 16352
rect 19376 16292 19380 16348
rect 19380 16292 19436 16348
rect 19436 16292 19440 16348
rect 19376 16288 19440 16292
rect 19456 16348 19520 16352
rect 19456 16292 19460 16348
rect 19460 16292 19516 16348
rect 19516 16292 19520 16348
rect 19456 16288 19520 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 10216 15804 10280 15808
rect 10216 15748 10220 15804
rect 10220 15748 10276 15804
rect 10276 15748 10280 15804
rect 10216 15744 10280 15748
rect 10296 15804 10360 15808
rect 10296 15748 10300 15804
rect 10300 15748 10356 15804
rect 10356 15748 10360 15804
rect 10296 15744 10360 15748
rect 10376 15804 10440 15808
rect 10376 15748 10380 15804
rect 10380 15748 10436 15804
rect 10436 15748 10440 15804
rect 10376 15744 10440 15748
rect 10456 15804 10520 15808
rect 10456 15748 10460 15804
rect 10460 15748 10516 15804
rect 10516 15748 10520 15804
rect 10456 15744 10520 15748
rect 16216 15804 16280 15808
rect 16216 15748 16220 15804
rect 16220 15748 16276 15804
rect 16276 15748 16280 15804
rect 16216 15744 16280 15748
rect 16296 15804 16360 15808
rect 16296 15748 16300 15804
rect 16300 15748 16356 15804
rect 16356 15748 16360 15804
rect 16296 15744 16360 15748
rect 16376 15804 16440 15808
rect 16376 15748 16380 15804
rect 16380 15748 16436 15804
rect 16436 15748 16440 15804
rect 16376 15744 16440 15748
rect 16456 15804 16520 15808
rect 16456 15748 16460 15804
rect 16460 15748 16516 15804
rect 16516 15748 16520 15804
rect 16456 15744 16520 15748
rect 7216 15260 7280 15264
rect 7216 15204 7220 15260
rect 7220 15204 7276 15260
rect 7276 15204 7280 15260
rect 7216 15200 7280 15204
rect 7296 15260 7360 15264
rect 7296 15204 7300 15260
rect 7300 15204 7356 15260
rect 7356 15204 7360 15260
rect 7296 15200 7360 15204
rect 7376 15260 7440 15264
rect 7376 15204 7380 15260
rect 7380 15204 7436 15260
rect 7436 15204 7440 15260
rect 7376 15200 7440 15204
rect 7456 15260 7520 15264
rect 7456 15204 7460 15260
rect 7460 15204 7516 15260
rect 7516 15204 7520 15260
rect 7456 15200 7520 15204
rect 13216 15260 13280 15264
rect 13216 15204 13220 15260
rect 13220 15204 13276 15260
rect 13276 15204 13280 15260
rect 13216 15200 13280 15204
rect 13296 15260 13360 15264
rect 13296 15204 13300 15260
rect 13300 15204 13356 15260
rect 13356 15204 13360 15260
rect 13296 15200 13360 15204
rect 13376 15260 13440 15264
rect 13376 15204 13380 15260
rect 13380 15204 13436 15260
rect 13436 15204 13440 15260
rect 13376 15200 13440 15204
rect 13456 15260 13520 15264
rect 13456 15204 13460 15260
rect 13460 15204 13516 15260
rect 13516 15204 13520 15260
rect 13456 15200 13520 15204
rect 19216 15260 19280 15264
rect 19216 15204 19220 15260
rect 19220 15204 19276 15260
rect 19276 15204 19280 15260
rect 19216 15200 19280 15204
rect 19296 15260 19360 15264
rect 19296 15204 19300 15260
rect 19300 15204 19356 15260
rect 19356 15204 19360 15260
rect 19296 15200 19360 15204
rect 19376 15260 19440 15264
rect 19376 15204 19380 15260
rect 19380 15204 19436 15260
rect 19436 15204 19440 15260
rect 19376 15200 19440 15204
rect 19456 15260 19520 15264
rect 19456 15204 19460 15260
rect 19460 15204 19516 15260
rect 19516 15204 19520 15260
rect 19456 15200 19520 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 10216 14716 10280 14720
rect 10216 14660 10220 14716
rect 10220 14660 10276 14716
rect 10276 14660 10280 14716
rect 10216 14656 10280 14660
rect 10296 14716 10360 14720
rect 10296 14660 10300 14716
rect 10300 14660 10356 14716
rect 10356 14660 10360 14716
rect 10296 14656 10360 14660
rect 10376 14716 10440 14720
rect 10376 14660 10380 14716
rect 10380 14660 10436 14716
rect 10436 14660 10440 14716
rect 10376 14656 10440 14660
rect 10456 14716 10520 14720
rect 10456 14660 10460 14716
rect 10460 14660 10516 14716
rect 10516 14660 10520 14716
rect 10456 14656 10520 14660
rect 16216 14716 16280 14720
rect 16216 14660 16220 14716
rect 16220 14660 16276 14716
rect 16276 14660 16280 14716
rect 16216 14656 16280 14660
rect 16296 14716 16360 14720
rect 16296 14660 16300 14716
rect 16300 14660 16356 14716
rect 16356 14660 16360 14716
rect 16296 14656 16360 14660
rect 16376 14716 16440 14720
rect 16376 14660 16380 14716
rect 16380 14660 16436 14716
rect 16436 14660 16440 14716
rect 16376 14656 16440 14660
rect 16456 14716 16520 14720
rect 16456 14660 16460 14716
rect 16460 14660 16516 14716
rect 16516 14660 16520 14716
rect 16456 14656 16520 14660
rect 7216 14172 7280 14176
rect 7216 14116 7220 14172
rect 7220 14116 7276 14172
rect 7276 14116 7280 14172
rect 7216 14112 7280 14116
rect 7296 14172 7360 14176
rect 7296 14116 7300 14172
rect 7300 14116 7356 14172
rect 7356 14116 7360 14172
rect 7296 14112 7360 14116
rect 7376 14172 7440 14176
rect 7376 14116 7380 14172
rect 7380 14116 7436 14172
rect 7436 14116 7440 14172
rect 7376 14112 7440 14116
rect 7456 14172 7520 14176
rect 7456 14116 7460 14172
rect 7460 14116 7516 14172
rect 7516 14116 7520 14172
rect 7456 14112 7520 14116
rect 13216 14172 13280 14176
rect 13216 14116 13220 14172
rect 13220 14116 13276 14172
rect 13276 14116 13280 14172
rect 13216 14112 13280 14116
rect 13296 14172 13360 14176
rect 13296 14116 13300 14172
rect 13300 14116 13356 14172
rect 13356 14116 13360 14172
rect 13296 14112 13360 14116
rect 13376 14172 13440 14176
rect 13376 14116 13380 14172
rect 13380 14116 13436 14172
rect 13436 14116 13440 14172
rect 13376 14112 13440 14116
rect 13456 14172 13520 14176
rect 13456 14116 13460 14172
rect 13460 14116 13516 14172
rect 13516 14116 13520 14172
rect 13456 14112 13520 14116
rect 19216 14172 19280 14176
rect 19216 14116 19220 14172
rect 19220 14116 19276 14172
rect 19276 14116 19280 14172
rect 19216 14112 19280 14116
rect 19296 14172 19360 14176
rect 19296 14116 19300 14172
rect 19300 14116 19356 14172
rect 19356 14116 19360 14172
rect 19296 14112 19360 14116
rect 19376 14172 19440 14176
rect 19376 14116 19380 14172
rect 19380 14116 19436 14172
rect 19436 14116 19440 14172
rect 19376 14112 19440 14116
rect 19456 14172 19520 14176
rect 19456 14116 19460 14172
rect 19460 14116 19516 14172
rect 19516 14116 19520 14172
rect 19456 14112 19520 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 10216 13628 10280 13632
rect 10216 13572 10220 13628
rect 10220 13572 10276 13628
rect 10276 13572 10280 13628
rect 10216 13568 10280 13572
rect 10296 13628 10360 13632
rect 10296 13572 10300 13628
rect 10300 13572 10356 13628
rect 10356 13572 10360 13628
rect 10296 13568 10360 13572
rect 10376 13628 10440 13632
rect 10376 13572 10380 13628
rect 10380 13572 10436 13628
rect 10436 13572 10440 13628
rect 10376 13568 10440 13572
rect 10456 13628 10520 13632
rect 10456 13572 10460 13628
rect 10460 13572 10516 13628
rect 10516 13572 10520 13628
rect 10456 13568 10520 13572
rect 16216 13628 16280 13632
rect 16216 13572 16220 13628
rect 16220 13572 16276 13628
rect 16276 13572 16280 13628
rect 16216 13568 16280 13572
rect 16296 13628 16360 13632
rect 16296 13572 16300 13628
rect 16300 13572 16356 13628
rect 16356 13572 16360 13628
rect 16296 13568 16360 13572
rect 16376 13628 16440 13632
rect 16376 13572 16380 13628
rect 16380 13572 16436 13628
rect 16436 13572 16440 13628
rect 16376 13568 16440 13572
rect 16456 13628 16520 13632
rect 16456 13572 16460 13628
rect 16460 13572 16516 13628
rect 16516 13572 16520 13628
rect 16456 13568 16520 13572
rect 7216 13084 7280 13088
rect 7216 13028 7220 13084
rect 7220 13028 7276 13084
rect 7276 13028 7280 13084
rect 7216 13024 7280 13028
rect 7296 13084 7360 13088
rect 7296 13028 7300 13084
rect 7300 13028 7356 13084
rect 7356 13028 7360 13084
rect 7296 13024 7360 13028
rect 7376 13084 7440 13088
rect 7376 13028 7380 13084
rect 7380 13028 7436 13084
rect 7436 13028 7440 13084
rect 7376 13024 7440 13028
rect 7456 13084 7520 13088
rect 7456 13028 7460 13084
rect 7460 13028 7516 13084
rect 7516 13028 7520 13084
rect 7456 13024 7520 13028
rect 13216 13084 13280 13088
rect 13216 13028 13220 13084
rect 13220 13028 13276 13084
rect 13276 13028 13280 13084
rect 13216 13024 13280 13028
rect 13296 13084 13360 13088
rect 13296 13028 13300 13084
rect 13300 13028 13356 13084
rect 13356 13028 13360 13084
rect 13296 13024 13360 13028
rect 13376 13084 13440 13088
rect 13376 13028 13380 13084
rect 13380 13028 13436 13084
rect 13436 13028 13440 13084
rect 13376 13024 13440 13028
rect 13456 13084 13520 13088
rect 13456 13028 13460 13084
rect 13460 13028 13516 13084
rect 13516 13028 13520 13084
rect 13456 13024 13520 13028
rect 19216 13084 19280 13088
rect 19216 13028 19220 13084
rect 19220 13028 19276 13084
rect 19276 13028 19280 13084
rect 19216 13024 19280 13028
rect 19296 13084 19360 13088
rect 19296 13028 19300 13084
rect 19300 13028 19356 13084
rect 19356 13028 19360 13084
rect 19296 13024 19360 13028
rect 19376 13084 19440 13088
rect 19376 13028 19380 13084
rect 19380 13028 19436 13084
rect 19436 13028 19440 13084
rect 19376 13024 19440 13028
rect 19456 13084 19520 13088
rect 19456 13028 19460 13084
rect 19460 13028 19516 13084
rect 19516 13028 19520 13084
rect 19456 13024 19520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 10216 12540 10280 12544
rect 10216 12484 10220 12540
rect 10220 12484 10276 12540
rect 10276 12484 10280 12540
rect 10216 12480 10280 12484
rect 10296 12540 10360 12544
rect 10296 12484 10300 12540
rect 10300 12484 10356 12540
rect 10356 12484 10360 12540
rect 10296 12480 10360 12484
rect 10376 12540 10440 12544
rect 10376 12484 10380 12540
rect 10380 12484 10436 12540
rect 10436 12484 10440 12540
rect 10376 12480 10440 12484
rect 10456 12540 10520 12544
rect 10456 12484 10460 12540
rect 10460 12484 10516 12540
rect 10516 12484 10520 12540
rect 10456 12480 10520 12484
rect 16216 12540 16280 12544
rect 16216 12484 16220 12540
rect 16220 12484 16276 12540
rect 16276 12484 16280 12540
rect 16216 12480 16280 12484
rect 16296 12540 16360 12544
rect 16296 12484 16300 12540
rect 16300 12484 16356 12540
rect 16356 12484 16360 12540
rect 16296 12480 16360 12484
rect 16376 12540 16440 12544
rect 16376 12484 16380 12540
rect 16380 12484 16436 12540
rect 16436 12484 16440 12540
rect 16376 12480 16440 12484
rect 16456 12540 16520 12544
rect 16456 12484 16460 12540
rect 16460 12484 16516 12540
rect 16516 12484 16520 12540
rect 16456 12480 16520 12484
rect 7216 11996 7280 12000
rect 7216 11940 7220 11996
rect 7220 11940 7276 11996
rect 7276 11940 7280 11996
rect 7216 11936 7280 11940
rect 7296 11996 7360 12000
rect 7296 11940 7300 11996
rect 7300 11940 7356 11996
rect 7356 11940 7360 11996
rect 7296 11936 7360 11940
rect 7376 11996 7440 12000
rect 7376 11940 7380 11996
rect 7380 11940 7436 11996
rect 7436 11940 7440 11996
rect 7376 11936 7440 11940
rect 7456 11996 7520 12000
rect 7456 11940 7460 11996
rect 7460 11940 7516 11996
rect 7516 11940 7520 11996
rect 7456 11936 7520 11940
rect 13216 11996 13280 12000
rect 13216 11940 13220 11996
rect 13220 11940 13276 11996
rect 13276 11940 13280 11996
rect 13216 11936 13280 11940
rect 13296 11996 13360 12000
rect 13296 11940 13300 11996
rect 13300 11940 13356 11996
rect 13356 11940 13360 11996
rect 13296 11936 13360 11940
rect 13376 11996 13440 12000
rect 13376 11940 13380 11996
rect 13380 11940 13436 11996
rect 13436 11940 13440 11996
rect 13376 11936 13440 11940
rect 13456 11996 13520 12000
rect 13456 11940 13460 11996
rect 13460 11940 13516 11996
rect 13516 11940 13520 11996
rect 13456 11936 13520 11940
rect 19216 11996 19280 12000
rect 19216 11940 19220 11996
rect 19220 11940 19276 11996
rect 19276 11940 19280 11996
rect 19216 11936 19280 11940
rect 19296 11996 19360 12000
rect 19296 11940 19300 11996
rect 19300 11940 19356 11996
rect 19356 11940 19360 11996
rect 19296 11936 19360 11940
rect 19376 11996 19440 12000
rect 19376 11940 19380 11996
rect 19380 11940 19436 11996
rect 19436 11940 19440 11996
rect 19376 11936 19440 11940
rect 19456 11996 19520 12000
rect 19456 11940 19460 11996
rect 19460 11940 19516 11996
rect 19516 11940 19520 11996
rect 19456 11936 19520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 10216 11452 10280 11456
rect 10216 11396 10220 11452
rect 10220 11396 10276 11452
rect 10276 11396 10280 11452
rect 10216 11392 10280 11396
rect 10296 11452 10360 11456
rect 10296 11396 10300 11452
rect 10300 11396 10356 11452
rect 10356 11396 10360 11452
rect 10296 11392 10360 11396
rect 10376 11452 10440 11456
rect 10376 11396 10380 11452
rect 10380 11396 10436 11452
rect 10436 11396 10440 11452
rect 10376 11392 10440 11396
rect 10456 11452 10520 11456
rect 10456 11396 10460 11452
rect 10460 11396 10516 11452
rect 10516 11396 10520 11452
rect 10456 11392 10520 11396
rect 16216 11452 16280 11456
rect 16216 11396 16220 11452
rect 16220 11396 16276 11452
rect 16276 11396 16280 11452
rect 16216 11392 16280 11396
rect 16296 11452 16360 11456
rect 16296 11396 16300 11452
rect 16300 11396 16356 11452
rect 16356 11396 16360 11452
rect 16296 11392 16360 11396
rect 16376 11452 16440 11456
rect 16376 11396 16380 11452
rect 16380 11396 16436 11452
rect 16436 11396 16440 11452
rect 16376 11392 16440 11396
rect 16456 11452 16520 11456
rect 16456 11396 16460 11452
rect 16460 11396 16516 11452
rect 16516 11396 16520 11452
rect 16456 11392 16520 11396
rect 7216 10908 7280 10912
rect 7216 10852 7220 10908
rect 7220 10852 7276 10908
rect 7276 10852 7280 10908
rect 7216 10848 7280 10852
rect 7296 10908 7360 10912
rect 7296 10852 7300 10908
rect 7300 10852 7356 10908
rect 7356 10852 7360 10908
rect 7296 10848 7360 10852
rect 7376 10908 7440 10912
rect 7376 10852 7380 10908
rect 7380 10852 7436 10908
rect 7436 10852 7440 10908
rect 7376 10848 7440 10852
rect 7456 10908 7520 10912
rect 7456 10852 7460 10908
rect 7460 10852 7516 10908
rect 7516 10852 7520 10908
rect 7456 10848 7520 10852
rect 13216 10908 13280 10912
rect 13216 10852 13220 10908
rect 13220 10852 13276 10908
rect 13276 10852 13280 10908
rect 13216 10848 13280 10852
rect 13296 10908 13360 10912
rect 13296 10852 13300 10908
rect 13300 10852 13356 10908
rect 13356 10852 13360 10908
rect 13296 10848 13360 10852
rect 13376 10908 13440 10912
rect 13376 10852 13380 10908
rect 13380 10852 13436 10908
rect 13436 10852 13440 10908
rect 13376 10848 13440 10852
rect 13456 10908 13520 10912
rect 13456 10852 13460 10908
rect 13460 10852 13516 10908
rect 13516 10852 13520 10908
rect 13456 10848 13520 10852
rect 19216 10908 19280 10912
rect 19216 10852 19220 10908
rect 19220 10852 19276 10908
rect 19276 10852 19280 10908
rect 19216 10848 19280 10852
rect 19296 10908 19360 10912
rect 19296 10852 19300 10908
rect 19300 10852 19356 10908
rect 19356 10852 19360 10908
rect 19296 10848 19360 10852
rect 19376 10908 19440 10912
rect 19376 10852 19380 10908
rect 19380 10852 19436 10908
rect 19436 10852 19440 10908
rect 19376 10848 19440 10852
rect 19456 10908 19520 10912
rect 19456 10852 19460 10908
rect 19460 10852 19516 10908
rect 19516 10852 19520 10908
rect 19456 10848 19520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 10216 10364 10280 10368
rect 10216 10308 10220 10364
rect 10220 10308 10276 10364
rect 10276 10308 10280 10364
rect 10216 10304 10280 10308
rect 10296 10364 10360 10368
rect 10296 10308 10300 10364
rect 10300 10308 10356 10364
rect 10356 10308 10360 10364
rect 10296 10304 10360 10308
rect 10376 10364 10440 10368
rect 10376 10308 10380 10364
rect 10380 10308 10436 10364
rect 10436 10308 10440 10364
rect 10376 10304 10440 10308
rect 10456 10364 10520 10368
rect 10456 10308 10460 10364
rect 10460 10308 10516 10364
rect 10516 10308 10520 10364
rect 10456 10304 10520 10308
rect 16216 10364 16280 10368
rect 16216 10308 16220 10364
rect 16220 10308 16276 10364
rect 16276 10308 16280 10364
rect 16216 10304 16280 10308
rect 16296 10364 16360 10368
rect 16296 10308 16300 10364
rect 16300 10308 16356 10364
rect 16356 10308 16360 10364
rect 16296 10304 16360 10308
rect 16376 10364 16440 10368
rect 16376 10308 16380 10364
rect 16380 10308 16436 10364
rect 16436 10308 16440 10364
rect 16376 10304 16440 10308
rect 16456 10364 16520 10368
rect 16456 10308 16460 10364
rect 16460 10308 16516 10364
rect 16516 10308 16520 10364
rect 16456 10304 16520 10308
rect 7216 9820 7280 9824
rect 7216 9764 7220 9820
rect 7220 9764 7276 9820
rect 7276 9764 7280 9820
rect 7216 9760 7280 9764
rect 7296 9820 7360 9824
rect 7296 9764 7300 9820
rect 7300 9764 7356 9820
rect 7356 9764 7360 9820
rect 7296 9760 7360 9764
rect 7376 9820 7440 9824
rect 7376 9764 7380 9820
rect 7380 9764 7436 9820
rect 7436 9764 7440 9820
rect 7376 9760 7440 9764
rect 7456 9820 7520 9824
rect 7456 9764 7460 9820
rect 7460 9764 7516 9820
rect 7516 9764 7520 9820
rect 7456 9760 7520 9764
rect 13216 9820 13280 9824
rect 13216 9764 13220 9820
rect 13220 9764 13276 9820
rect 13276 9764 13280 9820
rect 13216 9760 13280 9764
rect 13296 9820 13360 9824
rect 13296 9764 13300 9820
rect 13300 9764 13356 9820
rect 13356 9764 13360 9820
rect 13296 9760 13360 9764
rect 13376 9820 13440 9824
rect 13376 9764 13380 9820
rect 13380 9764 13436 9820
rect 13436 9764 13440 9820
rect 13376 9760 13440 9764
rect 13456 9820 13520 9824
rect 13456 9764 13460 9820
rect 13460 9764 13516 9820
rect 13516 9764 13520 9820
rect 13456 9760 13520 9764
rect 19216 9820 19280 9824
rect 19216 9764 19220 9820
rect 19220 9764 19276 9820
rect 19276 9764 19280 9820
rect 19216 9760 19280 9764
rect 19296 9820 19360 9824
rect 19296 9764 19300 9820
rect 19300 9764 19356 9820
rect 19356 9764 19360 9820
rect 19296 9760 19360 9764
rect 19376 9820 19440 9824
rect 19376 9764 19380 9820
rect 19380 9764 19436 9820
rect 19436 9764 19440 9820
rect 19376 9760 19440 9764
rect 19456 9820 19520 9824
rect 19456 9764 19460 9820
rect 19460 9764 19516 9820
rect 19516 9764 19520 9820
rect 19456 9760 19520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 10216 9276 10280 9280
rect 10216 9220 10220 9276
rect 10220 9220 10276 9276
rect 10276 9220 10280 9276
rect 10216 9216 10280 9220
rect 10296 9276 10360 9280
rect 10296 9220 10300 9276
rect 10300 9220 10356 9276
rect 10356 9220 10360 9276
rect 10296 9216 10360 9220
rect 10376 9276 10440 9280
rect 10376 9220 10380 9276
rect 10380 9220 10436 9276
rect 10436 9220 10440 9276
rect 10376 9216 10440 9220
rect 10456 9276 10520 9280
rect 10456 9220 10460 9276
rect 10460 9220 10516 9276
rect 10516 9220 10520 9276
rect 10456 9216 10520 9220
rect 16216 9276 16280 9280
rect 16216 9220 16220 9276
rect 16220 9220 16276 9276
rect 16276 9220 16280 9276
rect 16216 9216 16280 9220
rect 16296 9276 16360 9280
rect 16296 9220 16300 9276
rect 16300 9220 16356 9276
rect 16356 9220 16360 9276
rect 16296 9216 16360 9220
rect 16376 9276 16440 9280
rect 16376 9220 16380 9276
rect 16380 9220 16436 9276
rect 16436 9220 16440 9276
rect 16376 9216 16440 9220
rect 16456 9276 16520 9280
rect 16456 9220 16460 9276
rect 16460 9220 16516 9276
rect 16516 9220 16520 9276
rect 16456 9216 16520 9220
rect 7216 8732 7280 8736
rect 7216 8676 7220 8732
rect 7220 8676 7276 8732
rect 7276 8676 7280 8732
rect 7216 8672 7280 8676
rect 7296 8732 7360 8736
rect 7296 8676 7300 8732
rect 7300 8676 7356 8732
rect 7356 8676 7360 8732
rect 7296 8672 7360 8676
rect 7376 8732 7440 8736
rect 7376 8676 7380 8732
rect 7380 8676 7436 8732
rect 7436 8676 7440 8732
rect 7376 8672 7440 8676
rect 7456 8732 7520 8736
rect 7456 8676 7460 8732
rect 7460 8676 7516 8732
rect 7516 8676 7520 8732
rect 7456 8672 7520 8676
rect 13216 8732 13280 8736
rect 13216 8676 13220 8732
rect 13220 8676 13276 8732
rect 13276 8676 13280 8732
rect 13216 8672 13280 8676
rect 13296 8732 13360 8736
rect 13296 8676 13300 8732
rect 13300 8676 13356 8732
rect 13356 8676 13360 8732
rect 13296 8672 13360 8676
rect 13376 8732 13440 8736
rect 13376 8676 13380 8732
rect 13380 8676 13436 8732
rect 13436 8676 13440 8732
rect 13376 8672 13440 8676
rect 13456 8732 13520 8736
rect 13456 8676 13460 8732
rect 13460 8676 13516 8732
rect 13516 8676 13520 8732
rect 13456 8672 13520 8676
rect 19216 8732 19280 8736
rect 19216 8676 19220 8732
rect 19220 8676 19276 8732
rect 19276 8676 19280 8732
rect 19216 8672 19280 8676
rect 19296 8732 19360 8736
rect 19296 8676 19300 8732
rect 19300 8676 19356 8732
rect 19356 8676 19360 8732
rect 19296 8672 19360 8676
rect 19376 8732 19440 8736
rect 19376 8676 19380 8732
rect 19380 8676 19436 8732
rect 19436 8676 19440 8732
rect 19376 8672 19440 8676
rect 19456 8732 19520 8736
rect 19456 8676 19460 8732
rect 19460 8676 19516 8732
rect 19516 8676 19520 8732
rect 19456 8672 19520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 10216 8188 10280 8192
rect 10216 8132 10220 8188
rect 10220 8132 10276 8188
rect 10276 8132 10280 8188
rect 10216 8128 10280 8132
rect 10296 8188 10360 8192
rect 10296 8132 10300 8188
rect 10300 8132 10356 8188
rect 10356 8132 10360 8188
rect 10296 8128 10360 8132
rect 10376 8188 10440 8192
rect 10376 8132 10380 8188
rect 10380 8132 10436 8188
rect 10436 8132 10440 8188
rect 10376 8128 10440 8132
rect 10456 8188 10520 8192
rect 10456 8132 10460 8188
rect 10460 8132 10516 8188
rect 10516 8132 10520 8188
rect 10456 8128 10520 8132
rect 16216 8188 16280 8192
rect 16216 8132 16220 8188
rect 16220 8132 16276 8188
rect 16276 8132 16280 8188
rect 16216 8128 16280 8132
rect 16296 8188 16360 8192
rect 16296 8132 16300 8188
rect 16300 8132 16356 8188
rect 16356 8132 16360 8188
rect 16296 8128 16360 8132
rect 16376 8188 16440 8192
rect 16376 8132 16380 8188
rect 16380 8132 16436 8188
rect 16436 8132 16440 8188
rect 16376 8128 16440 8132
rect 16456 8188 16520 8192
rect 16456 8132 16460 8188
rect 16460 8132 16516 8188
rect 16516 8132 16520 8188
rect 16456 8128 16520 8132
rect 7216 7644 7280 7648
rect 7216 7588 7220 7644
rect 7220 7588 7276 7644
rect 7276 7588 7280 7644
rect 7216 7584 7280 7588
rect 7296 7644 7360 7648
rect 7296 7588 7300 7644
rect 7300 7588 7356 7644
rect 7356 7588 7360 7644
rect 7296 7584 7360 7588
rect 7376 7644 7440 7648
rect 7376 7588 7380 7644
rect 7380 7588 7436 7644
rect 7436 7588 7440 7644
rect 7376 7584 7440 7588
rect 7456 7644 7520 7648
rect 7456 7588 7460 7644
rect 7460 7588 7516 7644
rect 7516 7588 7520 7644
rect 7456 7584 7520 7588
rect 13216 7644 13280 7648
rect 13216 7588 13220 7644
rect 13220 7588 13276 7644
rect 13276 7588 13280 7644
rect 13216 7584 13280 7588
rect 13296 7644 13360 7648
rect 13296 7588 13300 7644
rect 13300 7588 13356 7644
rect 13356 7588 13360 7644
rect 13296 7584 13360 7588
rect 13376 7644 13440 7648
rect 13376 7588 13380 7644
rect 13380 7588 13436 7644
rect 13436 7588 13440 7644
rect 13376 7584 13440 7588
rect 13456 7644 13520 7648
rect 13456 7588 13460 7644
rect 13460 7588 13516 7644
rect 13516 7588 13520 7644
rect 13456 7584 13520 7588
rect 19216 7644 19280 7648
rect 19216 7588 19220 7644
rect 19220 7588 19276 7644
rect 19276 7588 19280 7644
rect 19216 7584 19280 7588
rect 19296 7644 19360 7648
rect 19296 7588 19300 7644
rect 19300 7588 19356 7644
rect 19356 7588 19360 7644
rect 19296 7584 19360 7588
rect 19376 7644 19440 7648
rect 19376 7588 19380 7644
rect 19380 7588 19436 7644
rect 19436 7588 19440 7644
rect 19376 7584 19440 7588
rect 19456 7644 19520 7648
rect 19456 7588 19460 7644
rect 19460 7588 19516 7644
rect 19516 7588 19520 7644
rect 19456 7584 19520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 10216 7100 10280 7104
rect 10216 7044 10220 7100
rect 10220 7044 10276 7100
rect 10276 7044 10280 7100
rect 10216 7040 10280 7044
rect 10296 7100 10360 7104
rect 10296 7044 10300 7100
rect 10300 7044 10356 7100
rect 10356 7044 10360 7100
rect 10296 7040 10360 7044
rect 10376 7100 10440 7104
rect 10376 7044 10380 7100
rect 10380 7044 10436 7100
rect 10436 7044 10440 7100
rect 10376 7040 10440 7044
rect 10456 7100 10520 7104
rect 10456 7044 10460 7100
rect 10460 7044 10516 7100
rect 10516 7044 10520 7100
rect 10456 7040 10520 7044
rect 16216 7100 16280 7104
rect 16216 7044 16220 7100
rect 16220 7044 16276 7100
rect 16276 7044 16280 7100
rect 16216 7040 16280 7044
rect 16296 7100 16360 7104
rect 16296 7044 16300 7100
rect 16300 7044 16356 7100
rect 16356 7044 16360 7100
rect 16296 7040 16360 7044
rect 16376 7100 16440 7104
rect 16376 7044 16380 7100
rect 16380 7044 16436 7100
rect 16436 7044 16440 7100
rect 16376 7040 16440 7044
rect 16456 7100 16520 7104
rect 16456 7044 16460 7100
rect 16460 7044 16516 7100
rect 16516 7044 16520 7100
rect 16456 7040 16520 7044
rect 7216 6556 7280 6560
rect 7216 6500 7220 6556
rect 7220 6500 7276 6556
rect 7276 6500 7280 6556
rect 7216 6496 7280 6500
rect 7296 6556 7360 6560
rect 7296 6500 7300 6556
rect 7300 6500 7356 6556
rect 7356 6500 7360 6556
rect 7296 6496 7360 6500
rect 7376 6556 7440 6560
rect 7376 6500 7380 6556
rect 7380 6500 7436 6556
rect 7436 6500 7440 6556
rect 7376 6496 7440 6500
rect 7456 6556 7520 6560
rect 7456 6500 7460 6556
rect 7460 6500 7516 6556
rect 7516 6500 7520 6556
rect 7456 6496 7520 6500
rect 13216 6556 13280 6560
rect 13216 6500 13220 6556
rect 13220 6500 13276 6556
rect 13276 6500 13280 6556
rect 13216 6496 13280 6500
rect 13296 6556 13360 6560
rect 13296 6500 13300 6556
rect 13300 6500 13356 6556
rect 13356 6500 13360 6556
rect 13296 6496 13360 6500
rect 13376 6556 13440 6560
rect 13376 6500 13380 6556
rect 13380 6500 13436 6556
rect 13436 6500 13440 6556
rect 13376 6496 13440 6500
rect 13456 6556 13520 6560
rect 13456 6500 13460 6556
rect 13460 6500 13516 6556
rect 13516 6500 13520 6556
rect 13456 6496 13520 6500
rect 19216 6556 19280 6560
rect 19216 6500 19220 6556
rect 19220 6500 19276 6556
rect 19276 6500 19280 6556
rect 19216 6496 19280 6500
rect 19296 6556 19360 6560
rect 19296 6500 19300 6556
rect 19300 6500 19356 6556
rect 19356 6500 19360 6556
rect 19296 6496 19360 6500
rect 19376 6556 19440 6560
rect 19376 6500 19380 6556
rect 19380 6500 19436 6556
rect 19436 6500 19440 6556
rect 19376 6496 19440 6500
rect 19456 6556 19520 6560
rect 19456 6500 19460 6556
rect 19460 6500 19516 6556
rect 19516 6500 19520 6556
rect 19456 6496 19520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 10216 6012 10280 6016
rect 10216 5956 10220 6012
rect 10220 5956 10276 6012
rect 10276 5956 10280 6012
rect 10216 5952 10280 5956
rect 10296 6012 10360 6016
rect 10296 5956 10300 6012
rect 10300 5956 10356 6012
rect 10356 5956 10360 6012
rect 10296 5952 10360 5956
rect 10376 6012 10440 6016
rect 10376 5956 10380 6012
rect 10380 5956 10436 6012
rect 10436 5956 10440 6012
rect 10376 5952 10440 5956
rect 10456 6012 10520 6016
rect 10456 5956 10460 6012
rect 10460 5956 10516 6012
rect 10516 5956 10520 6012
rect 10456 5952 10520 5956
rect 16216 6012 16280 6016
rect 16216 5956 16220 6012
rect 16220 5956 16276 6012
rect 16276 5956 16280 6012
rect 16216 5952 16280 5956
rect 16296 6012 16360 6016
rect 16296 5956 16300 6012
rect 16300 5956 16356 6012
rect 16356 5956 16360 6012
rect 16296 5952 16360 5956
rect 16376 6012 16440 6016
rect 16376 5956 16380 6012
rect 16380 5956 16436 6012
rect 16436 5956 16440 6012
rect 16376 5952 16440 5956
rect 16456 6012 16520 6016
rect 16456 5956 16460 6012
rect 16460 5956 16516 6012
rect 16516 5956 16520 6012
rect 16456 5952 16520 5956
rect 7216 5468 7280 5472
rect 7216 5412 7220 5468
rect 7220 5412 7276 5468
rect 7276 5412 7280 5468
rect 7216 5408 7280 5412
rect 7296 5468 7360 5472
rect 7296 5412 7300 5468
rect 7300 5412 7356 5468
rect 7356 5412 7360 5468
rect 7296 5408 7360 5412
rect 7376 5468 7440 5472
rect 7376 5412 7380 5468
rect 7380 5412 7436 5468
rect 7436 5412 7440 5468
rect 7376 5408 7440 5412
rect 7456 5468 7520 5472
rect 7456 5412 7460 5468
rect 7460 5412 7516 5468
rect 7516 5412 7520 5468
rect 7456 5408 7520 5412
rect 13216 5468 13280 5472
rect 13216 5412 13220 5468
rect 13220 5412 13276 5468
rect 13276 5412 13280 5468
rect 13216 5408 13280 5412
rect 13296 5468 13360 5472
rect 13296 5412 13300 5468
rect 13300 5412 13356 5468
rect 13356 5412 13360 5468
rect 13296 5408 13360 5412
rect 13376 5468 13440 5472
rect 13376 5412 13380 5468
rect 13380 5412 13436 5468
rect 13436 5412 13440 5468
rect 13376 5408 13440 5412
rect 13456 5468 13520 5472
rect 13456 5412 13460 5468
rect 13460 5412 13516 5468
rect 13516 5412 13520 5468
rect 13456 5408 13520 5412
rect 19216 5468 19280 5472
rect 19216 5412 19220 5468
rect 19220 5412 19276 5468
rect 19276 5412 19280 5468
rect 19216 5408 19280 5412
rect 19296 5468 19360 5472
rect 19296 5412 19300 5468
rect 19300 5412 19356 5468
rect 19356 5412 19360 5468
rect 19296 5408 19360 5412
rect 19376 5468 19440 5472
rect 19376 5412 19380 5468
rect 19380 5412 19436 5468
rect 19436 5412 19440 5468
rect 19376 5408 19440 5412
rect 19456 5468 19520 5472
rect 19456 5412 19460 5468
rect 19460 5412 19516 5468
rect 19516 5412 19520 5468
rect 19456 5408 19520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 10216 4924 10280 4928
rect 10216 4868 10220 4924
rect 10220 4868 10276 4924
rect 10276 4868 10280 4924
rect 10216 4864 10280 4868
rect 10296 4924 10360 4928
rect 10296 4868 10300 4924
rect 10300 4868 10356 4924
rect 10356 4868 10360 4924
rect 10296 4864 10360 4868
rect 10376 4924 10440 4928
rect 10376 4868 10380 4924
rect 10380 4868 10436 4924
rect 10436 4868 10440 4924
rect 10376 4864 10440 4868
rect 10456 4924 10520 4928
rect 10456 4868 10460 4924
rect 10460 4868 10516 4924
rect 10516 4868 10520 4924
rect 10456 4864 10520 4868
rect 16216 4924 16280 4928
rect 16216 4868 16220 4924
rect 16220 4868 16276 4924
rect 16276 4868 16280 4924
rect 16216 4864 16280 4868
rect 16296 4924 16360 4928
rect 16296 4868 16300 4924
rect 16300 4868 16356 4924
rect 16356 4868 16360 4924
rect 16296 4864 16360 4868
rect 16376 4924 16440 4928
rect 16376 4868 16380 4924
rect 16380 4868 16436 4924
rect 16436 4868 16440 4924
rect 16376 4864 16440 4868
rect 16456 4924 16520 4928
rect 16456 4868 16460 4924
rect 16460 4868 16516 4924
rect 16516 4868 16520 4924
rect 16456 4864 16520 4868
rect 7216 4380 7280 4384
rect 7216 4324 7220 4380
rect 7220 4324 7276 4380
rect 7276 4324 7280 4380
rect 7216 4320 7280 4324
rect 7296 4380 7360 4384
rect 7296 4324 7300 4380
rect 7300 4324 7356 4380
rect 7356 4324 7360 4380
rect 7296 4320 7360 4324
rect 7376 4380 7440 4384
rect 7376 4324 7380 4380
rect 7380 4324 7436 4380
rect 7436 4324 7440 4380
rect 7376 4320 7440 4324
rect 7456 4380 7520 4384
rect 7456 4324 7460 4380
rect 7460 4324 7516 4380
rect 7516 4324 7520 4380
rect 7456 4320 7520 4324
rect 13216 4380 13280 4384
rect 13216 4324 13220 4380
rect 13220 4324 13276 4380
rect 13276 4324 13280 4380
rect 13216 4320 13280 4324
rect 13296 4380 13360 4384
rect 13296 4324 13300 4380
rect 13300 4324 13356 4380
rect 13356 4324 13360 4380
rect 13296 4320 13360 4324
rect 13376 4380 13440 4384
rect 13376 4324 13380 4380
rect 13380 4324 13436 4380
rect 13436 4324 13440 4380
rect 13376 4320 13440 4324
rect 13456 4380 13520 4384
rect 13456 4324 13460 4380
rect 13460 4324 13516 4380
rect 13516 4324 13520 4380
rect 13456 4320 13520 4324
rect 19216 4380 19280 4384
rect 19216 4324 19220 4380
rect 19220 4324 19276 4380
rect 19276 4324 19280 4380
rect 19216 4320 19280 4324
rect 19296 4380 19360 4384
rect 19296 4324 19300 4380
rect 19300 4324 19356 4380
rect 19356 4324 19360 4380
rect 19296 4320 19360 4324
rect 19376 4380 19440 4384
rect 19376 4324 19380 4380
rect 19380 4324 19436 4380
rect 19436 4324 19440 4380
rect 19376 4320 19440 4324
rect 19456 4380 19520 4384
rect 19456 4324 19460 4380
rect 19460 4324 19516 4380
rect 19516 4324 19520 4380
rect 19456 4320 19520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 10216 3836 10280 3840
rect 10216 3780 10220 3836
rect 10220 3780 10276 3836
rect 10276 3780 10280 3836
rect 10216 3776 10280 3780
rect 10296 3836 10360 3840
rect 10296 3780 10300 3836
rect 10300 3780 10356 3836
rect 10356 3780 10360 3836
rect 10296 3776 10360 3780
rect 10376 3836 10440 3840
rect 10376 3780 10380 3836
rect 10380 3780 10436 3836
rect 10436 3780 10440 3836
rect 10376 3776 10440 3780
rect 10456 3836 10520 3840
rect 10456 3780 10460 3836
rect 10460 3780 10516 3836
rect 10516 3780 10520 3836
rect 10456 3776 10520 3780
rect 16216 3836 16280 3840
rect 16216 3780 16220 3836
rect 16220 3780 16276 3836
rect 16276 3780 16280 3836
rect 16216 3776 16280 3780
rect 16296 3836 16360 3840
rect 16296 3780 16300 3836
rect 16300 3780 16356 3836
rect 16356 3780 16360 3836
rect 16296 3776 16360 3780
rect 16376 3836 16440 3840
rect 16376 3780 16380 3836
rect 16380 3780 16436 3836
rect 16436 3780 16440 3836
rect 16376 3776 16440 3780
rect 16456 3836 16520 3840
rect 16456 3780 16460 3836
rect 16460 3780 16516 3836
rect 16516 3780 16520 3836
rect 16456 3776 16520 3780
rect 7216 3292 7280 3296
rect 7216 3236 7220 3292
rect 7220 3236 7276 3292
rect 7276 3236 7280 3292
rect 7216 3232 7280 3236
rect 7296 3292 7360 3296
rect 7296 3236 7300 3292
rect 7300 3236 7356 3292
rect 7356 3236 7360 3292
rect 7296 3232 7360 3236
rect 7376 3292 7440 3296
rect 7376 3236 7380 3292
rect 7380 3236 7436 3292
rect 7436 3236 7440 3292
rect 7376 3232 7440 3236
rect 7456 3292 7520 3296
rect 7456 3236 7460 3292
rect 7460 3236 7516 3292
rect 7516 3236 7520 3292
rect 7456 3232 7520 3236
rect 13216 3292 13280 3296
rect 13216 3236 13220 3292
rect 13220 3236 13276 3292
rect 13276 3236 13280 3292
rect 13216 3232 13280 3236
rect 13296 3292 13360 3296
rect 13296 3236 13300 3292
rect 13300 3236 13356 3292
rect 13356 3236 13360 3292
rect 13296 3232 13360 3236
rect 13376 3292 13440 3296
rect 13376 3236 13380 3292
rect 13380 3236 13436 3292
rect 13436 3236 13440 3292
rect 13376 3232 13440 3236
rect 13456 3292 13520 3296
rect 13456 3236 13460 3292
rect 13460 3236 13516 3292
rect 13516 3236 13520 3292
rect 13456 3232 13520 3236
rect 19216 3292 19280 3296
rect 19216 3236 19220 3292
rect 19220 3236 19276 3292
rect 19276 3236 19280 3292
rect 19216 3232 19280 3236
rect 19296 3292 19360 3296
rect 19296 3236 19300 3292
rect 19300 3236 19356 3292
rect 19356 3236 19360 3292
rect 19296 3232 19360 3236
rect 19376 3292 19440 3296
rect 19376 3236 19380 3292
rect 19380 3236 19436 3292
rect 19436 3236 19440 3292
rect 19376 3232 19440 3236
rect 19456 3292 19520 3296
rect 19456 3236 19460 3292
rect 19460 3236 19516 3292
rect 19516 3236 19520 3292
rect 19456 3232 19520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 10216 2748 10280 2752
rect 10216 2692 10220 2748
rect 10220 2692 10276 2748
rect 10276 2692 10280 2748
rect 10216 2688 10280 2692
rect 10296 2748 10360 2752
rect 10296 2692 10300 2748
rect 10300 2692 10356 2748
rect 10356 2692 10360 2748
rect 10296 2688 10360 2692
rect 10376 2748 10440 2752
rect 10376 2692 10380 2748
rect 10380 2692 10436 2748
rect 10436 2692 10440 2748
rect 10376 2688 10440 2692
rect 10456 2748 10520 2752
rect 10456 2692 10460 2748
rect 10460 2692 10516 2748
rect 10516 2692 10520 2748
rect 10456 2688 10520 2692
rect 16216 2748 16280 2752
rect 16216 2692 16220 2748
rect 16220 2692 16276 2748
rect 16276 2692 16280 2748
rect 16216 2688 16280 2692
rect 16296 2748 16360 2752
rect 16296 2692 16300 2748
rect 16300 2692 16356 2748
rect 16356 2692 16360 2748
rect 16296 2688 16360 2692
rect 16376 2748 16440 2752
rect 16376 2692 16380 2748
rect 16380 2692 16436 2748
rect 16436 2692 16440 2748
rect 16376 2688 16440 2692
rect 16456 2748 16520 2752
rect 16456 2692 16460 2748
rect 16460 2692 16516 2748
rect 16516 2692 16520 2748
rect 16456 2688 16520 2692
rect 7216 2204 7280 2208
rect 7216 2148 7220 2204
rect 7220 2148 7276 2204
rect 7276 2148 7280 2204
rect 7216 2144 7280 2148
rect 7296 2204 7360 2208
rect 7296 2148 7300 2204
rect 7300 2148 7356 2204
rect 7356 2148 7360 2204
rect 7296 2144 7360 2148
rect 7376 2204 7440 2208
rect 7376 2148 7380 2204
rect 7380 2148 7436 2204
rect 7436 2148 7440 2204
rect 7376 2144 7440 2148
rect 7456 2204 7520 2208
rect 7456 2148 7460 2204
rect 7460 2148 7516 2204
rect 7516 2148 7520 2204
rect 7456 2144 7520 2148
rect 13216 2204 13280 2208
rect 13216 2148 13220 2204
rect 13220 2148 13276 2204
rect 13276 2148 13280 2204
rect 13216 2144 13280 2148
rect 13296 2204 13360 2208
rect 13296 2148 13300 2204
rect 13300 2148 13356 2204
rect 13356 2148 13360 2204
rect 13296 2144 13360 2148
rect 13376 2204 13440 2208
rect 13376 2148 13380 2204
rect 13380 2148 13436 2204
rect 13436 2148 13440 2204
rect 13376 2144 13440 2148
rect 13456 2204 13520 2208
rect 13456 2148 13460 2204
rect 13460 2148 13516 2204
rect 13516 2148 13520 2204
rect 13456 2144 13520 2148
rect 19216 2204 19280 2208
rect 19216 2148 19220 2204
rect 19220 2148 19276 2204
rect 19276 2148 19280 2204
rect 19216 2144 19280 2148
rect 19296 2204 19360 2208
rect 19296 2148 19300 2204
rect 19300 2148 19356 2204
rect 19356 2148 19360 2204
rect 19296 2144 19360 2148
rect 19376 2204 19440 2208
rect 19376 2148 19380 2204
rect 19380 2148 19436 2204
rect 19436 2148 19440 2204
rect 19376 2144 19440 2148
rect 19456 2204 19520 2208
rect 19456 2148 19460 2204
rect 19460 2148 19516 2204
rect 19516 2148 19520 2204
rect 19456 2144 19520 2148
<< metal4 >>
rect 4208 21248 4528 21808
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 7208 21792 7528 21808
rect 7208 21728 7216 21792
rect 7280 21728 7296 21792
rect 7360 21728 7376 21792
rect 7440 21728 7456 21792
rect 7520 21728 7528 21792
rect 7208 20704 7528 21728
rect 7208 20640 7216 20704
rect 7280 20640 7296 20704
rect 7360 20640 7376 20704
rect 7440 20640 7456 20704
rect 7520 20640 7528 20704
rect 7208 19616 7528 20640
rect 7208 19552 7216 19616
rect 7280 19552 7296 19616
rect 7360 19552 7376 19616
rect 7440 19552 7456 19616
rect 7520 19552 7528 19616
rect 7208 18528 7528 19552
rect 7208 18464 7216 18528
rect 7280 18464 7296 18528
rect 7360 18464 7376 18528
rect 7440 18464 7456 18528
rect 7520 18464 7528 18528
rect 7208 17440 7528 18464
rect 7208 17376 7216 17440
rect 7280 17376 7296 17440
rect 7360 17376 7376 17440
rect 7440 17376 7456 17440
rect 7520 17376 7528 17440
rect 7208 16352 7528 17376
rect 7208 16288 7216 16352
rect 7280 16288 7296 16352
rect 7360 16288 7376 16352
rect 7440 16288 7456 16352
rect 7520 16288 7528 16352
rect 7208 15264 7528 16288
rect 7208 15200 7216 15264
rect 7280 15200 7296 15264
rect 7360 15200 7376 15264
rect 7440 15200 7456 15264
rect 7520 15200 7528 15264
rect 7208 14176 7528 15200
rect 7208 14112 7216 14176
rect 7280 14112 7296 14176
rect 7360 14112 7376 14176
rect 7440 14112 7456 14176
rect 7520 14112 7528 14176
rect 7208 13088 7528 14112
rect 7208 13024 7216 13088
rect 7280 13024 7296 13088
rect 7360 13024 7376 13088
rect 7440 13024 7456 13088
rect 7520 13024 7528 13088
rect 7208 12000 7528 13024
rect 7208 11936 7216 12000
rect 7280 11936 7296 12000
rect 7360 11936 7376 12000
rect 7440 11936 7456 12000
rect 7520 11936 7528 12000
rect 7208 10912 7528 11936
rect 7208 10848 7216 10912
rect 7280 10848 7296 10912
rect 7360 10848 7376 10912
rect 7440 10848 7456 10912
rect 7520 10848 7528 10912
rect 7208 9824 7528 10848
rect 7208 9760 7216 9824
rect 7280 9760 7296 9824
rect 7360 9760 7376 9824
rect 7440 9760 7456 9824
rect 7520 9760 7528 9824
rect 7208 8736 7528 9760
rect 7208 8672 7216 8736
rect 7280 8672 7296 8736
rect 7360 8672 7376 8736
rect 7440 8672 7456 8736
rect 7520 8672 7528 8736
rect 7208 7648 7528 8672
rect 7208 7584 7216 7648
rect 7280 7584 7296 7648
rect 7360 7584 7376 7648
rect 7440 7584 7456 7648
rect 7520 7584 7528 7648
rect 7208 6560 7528 7584
rect 7208 6496 7216 6560
rect 7280 6496 7296 6560
rect 7360 6496 7376 6560
rect 7440 6496 7456 6560
rect 7520 6496 7528 6560
rect 7208 5472 7528 6496
rect 7208 5408 7216 5472
rect 7280 5408 7296 5472
rect 7360 5408 7376 5472
rect 7440 5408 7456 5472
rect 7520 5408 7528 5472
rect 7208 4384 7528 5408
rect 7208 4320 7216 4384
rect 7280 4320 7296 4384
rect 7360 4320 7376 4384
rect 7440 4320 7456 4384
rect 7520 4320 7528 4384
rect 7208 3296 7528 4320
rect 7208 3232 7216 3296
rect 7280 3232 7296 3296
rect 7360 3232 7376 3296
rect 7440 3232 7456 3296
rect 7520 3232 7528 3296
rect 7208 2208 7528 3232
rect 7208 2144 7216 2208
rect 7280 2144 7296 2208
rect 7360 2144 7376 2208
rect 7440 2144 7456 2208
rect 7520 2144 7528 2208
rect 7208 2128 7528 2144
rect 10208 21248 10528 21808
rect 10208 21184 10216 21248
rect 10280 21184 10296 21248
rect 10360 21184 10376 21248
rect 10440 21184 10456 21248
rect 10520 21184 10528 21248
rect 10208 20160 10528 21184
rect 10208 20096 10216 20160
rect 10280 20096 10296 20160
rect 10360 20096 10376 20160
rect 10440 20096 10456 20160
rect 10520 20096 10528 20160
rect 10208 19072 10528 20096
rect 10208 19008 10216 19072
rect 10280 19008 10296 19072
rect 10360 19008 10376 19072
rect 10440 19008 10456 19072
rect 10520 19008 10528 19072
rect 10208 17984 10528 19008
rect 10208 17920 10216 17984
rect 10280 17920 10296 17984
rect 10360 17920 10376 17984
rect 10440 17920 10456 17984
rect 10520 17920 10528 17984
rect 10208 16896 10528 17920
rect 10208 16832 10216 16896
rect 10280 16832 10296 16896
rect 10360 16832 10376 16896
rect 10440 16832 10456 16896
rect 10520 16832 10528 16896
rect 10208 15808 10528 16832
rect 10208 15744 10216 15808
rect 10280 15744 10296 15808
rect 10360 15744 10376 15808
rect 10440 15744 10456 15808
rect 10520 15744 10528 15808
rect 10208 14720 10528 15744
rect 10208 14656 10216 14720
rect 10280 14656 10296 14720
rect 10360 14656 10376 14720
rect 10440 14656 10456 14720
rect 10520 14656 10528 14720
rect 10208 13632 10528 14656
rect 10208 13568 10216 13632
rect 10280 13568 10296 13632
rect 10360 13568 10376 13632
rect 10440 13568 10456 13632
rect 10520 13568 10528 13632
rect 10208 12544 10528 13568
rect 10208 12480 10216 12544
rect 10280 12480 10296 12544
rect 10360 12480 10376 12544
rect 10440 12480 10456 12544
rect 10520 12480 10528 12544
rect 10208 11456 10528 12480
rect 10208 11392 10216 11456
rect 10280 11392 10296 11456
rect 10360 11392 10376 11456
rect 10440 11392 10456 11456
rect 10520 11392 10528 11456
rect 10208 10368 10528 11392
rect 10208 10304 10216 10368
rect 10280 10304 10296 10368
rect 10360 10304 10376 10368
rect 10440 10304 10456 10368
rect 10520 10304 10528 10368
rect 10208 9280 10528 10304
rect 10208 9216 10216 9280
rect 10280 9216 10296 9280
rect 10360 9216 10376 9280
rect 10440 9216 10456 9280
rect 10520 9216 10528 9280
rect 10208 8192 10528 9216
rect 10208 8128 10216 8192
rect 10280 8128 10296 8192
rect 10360 8128 10376 8192
rect 10440 8128 10456 8192
rect 10520 8128 10528 8192
rect 10208 7104 10528 8128
rect 10208 7040 10216 7104
rect 10280 7040 10296 7104
rect 10360 7040 10376 7104
rect 10440 7040 10456 7104
rect 10520 7040 10528 7104
rect 10208 6016 10528 7040
rect 10208 5952 10216 6016
rect 10280 5952 10296 6016
rect 10360 5952 10376 6016
rect 10440 5952 10456 6016
rect 10520 5952 10528 6016
rect 10208 4928 10528 5952
rect 10208 4864 10216 4928
rect 10280 4864 10296 4928
rect 10360 4864 10376 4928
rect 10440 4864 10456 4928
rect 10520 4864 10528 4928
rect 10208 3840 10528 4864
rect 10208 3776 10216 3840
rect 10280 3776 10296 3840
rect 10360 3776 10376 3840
rect 10440 3776 10456 3840
rect 10520 3776 10528 3840
rect 10208 2752 10528 3776
rect 10208 2688 10216 2752
rect 10280 2688 10296 2752
rect 10360 2688 10376 2752
rect 10440 2688 10456 2752
rect 10520 2688 10528 2752
rect 10208 2128 10528 2688
rect 13208 21792 13528 21808
rect 13208 21728 13216 21792
rect 13280 21728 13296 21792
rect 13360 21728 13376 21792
rect 13440 21728 13456 21792
rect 13520 21728 13528 21792
rect 13208 20704 13528 21728
rect 13208 20640 13216 20704
rect 13280 20640 13296 20704
rect 13360 20640 13376 20704
rect 13440 20640 13456 20704
rect 13520 20640 13528 20704
rect 13208 19616 13528 20640
rect 13208 19552 13216 19616
rect 13280 19552 13296 19616
rect 13360 19552 13376 19616
rect 13440 19552 13456 19616
rect 13520 19552 13528 19616
rect 13208 18528 13528 19552
rect 13208 18464 13216 18528
rect 13280 18464 13296 18528
rect 13360 18464 13376 18528
rect 13440 18464 13456 18528
rect 13520 18464 13528 18528
rect 13208 17440 13528 18464
rect 13208 17376 13216 17440
rect 13280 17376 13296 17440
rect 13360 17376 13376 17440
rect 13440 17376 13456 17440
rect 13520 17376 13528 17440
rect 13208 16352 13528 17376
rect 13208 16288 13216 16352
rect 13280 16288 13296 16352
rect 13360 16288 13376 16352
rect 13440 16288 13456 16352
rect 13520 16288 13528 16352
rect 13208 15264 13528 16288
rect 13208 15200 13216 15264
rect 13280 15200 13296 15264
rect 13360 15200 13376 15264
rect 13440 15200 13456 15264
rect 13520 15200 13528 15264
rect 13208 14176 13528 15200
rect 13208 14112 13216 14176
rect 13280 14112 13296 14176
rect 13360 14112 13376 14176
rect 13440 14112 13456 14176
rect 13520 14112 13528 14176
rect 13208 13088 13528 14112
rect 13208 13024 13216 13088
rect 13280 13024 13296 13088
rect 13360 13024 13376 13088
rect 13440 13024 13456 13088
rect 13520 13024 13528 13088
rect 13208 12000 13528 13024
rect 13208 11936 13216 12000
rect 13280 11936 13296 12000
rect 13360 11936 13376 12000
rect 13440 11936 13456 12000
rect 13520 11936 13528 12000
rect 13208 10912 13528 11936
rect 13208 10848 13216 10912
rect 13280 10848 13296 10912
rect 13360 10848 13376 10912
rect 13440 10848 13456 10912
rect 13520 10848 13528 10912
rect 13208 9824 13528 10848
rect 13208 9760 13216 9824
rect 13280 9760 13296 9824
rect 13360 9760 13376 9824
rect 13440 9760 13456 9824
rect 13520 9760 13528 9824
rect 13208 8736 13528 9760
rect 13208 8672 13216 8736
rect 13280 8672 13296 8736
rect 13360 8672 13376 8736
rect 13440 8672 13456 8736
rect 13520 8672 13528 8736
rect 13208 7648 13528 8672
rect 13208 7584 13216 7648
rect 13280 7584 13296 7648
rect 13360 7584 13376 7648
rect 13440 7584 13456 7648
rect 13520 7584 13528 7648
rect 13208 6560 13528 7584
rect 13208 6496 13216 6560
rect 13280 6496 13296 6560
rect 13360 6496 13376 6560
rect 13440 6496 13456 6560
rect 13520 6496 13528 6560
rect 13208 5472 13528 6496
rect 13208 5408 13216 5472
rect 13280 5408 13296 5472
rect 13360 5408 13376 5472
rect 13440 5408 13456 5472
rect 13520 5408 13528 5472
rect 13208 4384 13528 5408
rect 13208 4320 13216 4384
rect 13280 4320 13296 4384
rect 13360 4320 13376 4384
rect 13440 4320 13456 4384
rect 13520 4320 13528 4384
rect 13208 3296 13528 4320
rect 13208 3232 13216 3296
rect 13280 3232 13296 3296
rect 13360 3232 13376 3296
rect 13440 3232 13456 3296
rect 13520 3232 13528 3296
rect 13208 2208 13528 3232
rect 13208 2144 13216 2208
rect 13280 2144 13296 2208
rect 13360 2144 13376 2208
rect 13440 2144 13456 2208
rect 13520 2144 13528 2208
rect 13208 2128 13528 2144
rect 16208 21248 16528 21808
rect 16208 21184 16216 21248
rect 16280 21184 16296 21248
rect 16360 21184 16376 21248
rect 16440 21184 16456 21248
rect 16520 21184 16528 21248
rect 16208 20160 16528 21184
rect 16208 20096 16216 20160
rect 16280 20096 16296 20160
rect 16360 20096 16376 20160
rect 16440 20096 16456 20160
rect 16520 20096 16528 20160
rect 16208 19072 16528 20096
rect 16208 19008 16216 19072
rect 16280 19008 16296 19072
rect 16360 19008 16376 19072
rect 16440 19008 16456 19072
rect 16520 19008 16528 19072
rect 16208 17984 16528 19008
rect 16208 17920 16216 17984
rect 16280 17920 16296 17984
rect 16360 17920 16376 17984
rect 16440 17920 16456 17984
rect 16520 17920 16528 17984
rect 16208 16896 16528 17920
rect 16208 16832 16216 16896
rect 16280 16832 16296 16896
rect 16360 16832 16376 16896
rect 16440 16832 16456 16896
rect 16520 16832 16528 16896
rect 16208 15808 16528 16832
rect 16208 15744 16216 15808
rect 16280 15744 16296 15808
rect 16360 15744 16376 15808
rect 16440 15744 16456 15808
rect 16520 15744 16528 15808
rect 16208 14720 16528 15744
rect 16208 14656 16216 14720
rect 16280 14656 16296 14720
rect 16360 14656 16376 14720
rect 16440 14656 16456 14720
rect 16520 14656 16528 14720
rect 16208 13632 16528 14656
rect 16208 13568 16216 13632
rect 16280 13568 16296 13632
rect 16360 13568 16376 13632
rect 16440 13568 16456 13632
rect 16520 13568 16528 13632
rect 16208 12544 16528 13568
rect 16208 12480 16216 12544
rect 16280 12480 16296 12544
rect 16360 12480 16376 12544
rect 16440 12480 16456 12544
rect 16520 12480 16528 12544
rect 16208 11456 16528 12480
rect 16208 11392 16216 11456
rect 16280 11392 16296 11456
rect 16360 11392 16376 11456
rect 16440 11392 16456 11456
rect 16520 11392 16528 11456
rect 16208 10368 16528 11392
rect 16208 10304 16216 10368
rect 16280 10304 16296 10368
rect 16360 10304 16376 10368
rect 16440 10304 16456 10368
rect 16520 10304 16528 10368
rect 16208 9280 16528 10304
rect 16208 9216 16216 9280
rect 16280 9216 16296 9280
rect 16360 9216 16376 9280
rect 16440 9216 16456 9280
rect 16520 9216 16528 9280
rect 16208 8192 16528 9216
rect 16208 8128 16216 8192
rect 16280 8128 16296 8192
rect 16360 8128 16376 8192
rect 16440 8128 16456 8192
rect 16520 8128 16528 8192
rect 16208 7104 16528 8128
rect 16208 7040 16216 7104
rect 16280 7040 16296 7104
rect 16360 7040 16376 7104
rect 16440 7040 16456 7104
rect 16520 7040 16528 7104
rect 16208 6016 16528 7040
rect 16208 5952 16216 6016
rect 16280 5952 16296 6016
rect 16360 5952 16376 6016
rect 16440 5952 16456 6016
rect 16520 5952 16528 6016
rect 16208 4928 16528 5952
rect 16208 4864 16216 4928
rect 16280 4864 16296 4928
rect 16360 4864 16376 4928
rect 16440 4864 16456 4928
rect 16520 4864 16528 4928
rect 16208 3840 16528 4864
rect 16208 3776 16216 3840
rect 16280 3776 16296 3840
rect 16360 3776 16376 3840
rect 16440 3776 16456 3840
rect 16520 3776 16528 3840
rect 16208 2752 16528 3776
rect 16208 2688 16216 2752
rect 16280 2688 16296 2752
rect 16360 2688 16376 2752
rect 16440 2688 16456 2752
rect 16520 2688 16528 2752
rect 16208 2128 16528 2688
rect 19208 21792 19528 21808
rect 19208 21728 19216 21792
rect 19280 21728 19296 21792
rect 19360 21728 19376 21792
rect 19440 21728 19456 21792
rect 19520 21728 19528 21792
rect 19208 20704 19528 21728
rect 19208 20640 19216 20704
rect 19280 20640 19296 20704
rect 19360 20640 19376 20704
rect 19440 20640 19456 20704
rect 19520 20640 19528 20704
rect 19208 19616 19528 20640
rect 19208 19552 19216 19616
rect 19280 19552 19296 19616
rect 19360 19552 19376 19616
rect 19440 19552 19456 19616
rect 19520 19552 19528 19616
rect 19208 18528 19528 19552
rect 19208 18464 19216 18528
rect 19280 18464 19296 18528
rect 19360 18464 19376 18528
rect 19440 18464 19456 18528
rect 19520 18464 19528 18528
rect 19208 17440 19528 18464
rect 19208 17376 19216 17440
rect 19280 17376 19296 17440
rect 19360 17376 19376 17440
rect 19440 17376 19456 17440
rect 19520 17376 19528 17440
rect 19208 16352 19528 17376
rect 19208 16288 19216 16352
rect 19280 16288 19296 16352
rect 19360 16288 19376 16352
rect 19440 16288 19456 16352
rect 19520 16288 19528 16352
rect 19208 15264 19528 16288
rect 19208 15200 19216 15264
rect 19280 15200 19296 15264
rect 19360 15200 19376 15264
rect 19440 15200 19456 15264
rect 19520 15200 19528 15264
rect 19208 14176 19528 15200
rect 19208 14112 19216 14176
rect 19280 14112 19296 14176
rect 19360 14112 19376 14176
rect 19440 14112 19456 14176
rect 19520 14112 19528 14176
rect 19208 13088 19528 14112
rect 19208 13024 19216 13088
rect 19280 13024 19296 13088
rect 19360 13024 19376 13088
rect 19440 13024 19456 13088
rect 19520 13024 19528 13088
rect 19208 12000 19528 13024
rect 19208 11936 19216 12000
rect 19280 11936 19296 12000
rect 19360 11936 19376 12000
rect 19440 11936 19456 12000
rect 19520 11936 19528 12000
rect 19208 10912 19528 11936
rect 19208 10848 19216 10912
rect 19280 10848 19296 10912
rect 19360 10848 19376 10912
rect 19440 10848 19456 10912
rect 19520 10848 19528 10912
rect 19208 9824 19528 10848
rect 19208 9760 19216 9824
rect 19280 9760 19296 9824
rect 19360 9760 19376 9824
rect 19440 9760 19456 9824
rect 19520 9760 19528 9824
rect 19208 8736 19528 9760
rect 19208 8672 19216 8736
rect 19280 8672 19296 8736
rect 19360 8672 19376 8736
rect 19440 8672 19456 8736
rect 19520 8672 19528 8736
rect 19208 7648 19528 8672
rect 19208 7584 19216 7648
rect 19280 7584 19296 7648
rect 19360 7584 19376 7648
rect 19440 7584 19456 7648
rect 19520 7584 19528 7648
rect 19208 6560 19528 7584
rect 19208 6496 19216 6560
rect 19280 6496 19296 6560
rect 19360 6496 19376 6560
rect 19440 6496 19456 6560
rect 19520 6496 19528 6560
rect 19208 5472 19528 6496
rect 19208 5408 19216 5472
rect 19280 5408 19296 5472
rect 19360 5408 19376 5472
rect 19440 5408 19456 5472
rect 19520 5408 19528 5472
rect 19208 4384 19528 5408
rect 19208 4320 19216 4384
rect 19280 4320 19296 4384
rect 19360 4320 19376 4384
rect 19440 4320 19456 4384
rect 19520 4320 19528 4384
rect 19208 3296 19528 4320
rect 19208 3232 19216 3296
rect 19280 3232 19296 3296
rect 19360 3232 19376 3296
rect 19440 3232 19456 3296
rect 19520 3232 19528 3296
rect 19208 2208 19528 3232
rect 19208 2144 19216 2208
rect 19280 2144 19296 2208
rect 19360 2144 19376 2208
rect 19440 2144 19456 2208
rect 19520 2144 19528 2208
rect 19208 2128 19528 2144
use sky130_fd_sc_hd__and4_1  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 18952 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 15824 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _169_
timestamp 1693170804
transform -1 0 13984 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _170_
timestamp 1693170804
transform -1 0 16560 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1693170804
transform 1 0 16652 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18124 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _174_
timestamp 1693170804
transform 1 0 15640 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _175_
timestamp 1693170804
transform 1 0 16836 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _176_
timestamp 1693170804
transform 1 0 17112 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 19780 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 17848 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _179_
timestamp 1693170804
transform -1 0 16284 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _180_
timestamp 1693170804
transform -1 0 13800 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _181_
timestamp 1693170804
transform 1 0 13064 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _182_
timestamp 1693170804
transform 1 0 12788 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _183_
timestamp 1693170804
transform 1 0 13248 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _184_
timestamp 1693170804
transform 1 0 14444 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _185_
timestamp 1693170804
transform 1 0 14076 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _186_
timestamp 1693170804
transform 1 0 12604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _187_
timestamp 1693170804
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _188_
timestamp 1693170804
transform 1 0 13708 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _189_
timestamp 1693170804
transform 1 0 14904 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _190_
timestamp 1693170804
transform -1 0 16192 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _191_
timestamp 1693170804
transform 1 0 19780 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _192_
timestamp 1693170804
transform 1 0 16008 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _193_
timestamp 1693170804
transform 1 0 16744 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _194_
timestamp 1693170804
transform -1 0 19872 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _195_
timestamp 1693170804
transform 1 0 18032 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _196_
timestamp 1693170804
transform -1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _197_
timestamp 1693170804
transform 1 0 16652 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _198_
timestamp 1693170804
transform 1 0 16744 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _199_
timestamp 1693170804
transform 1 0 19872 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _200_
timestamp 1693170804
transform 1 0 17112 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _201_
timestamp 1693170804
transform 1 0 17572 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _202_
timestamp 1693170804
transform 1 0 18308 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _203_
timestamp 1693170804
transform -1 0 19872 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _204_
timestamp 1693170804
transform -1 0 18124 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _205_
timestamp 1693170804
transform 1 0 16928 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _206_
timestamp 1693170804
transform -1 0 20332 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _207_
timestamp 1693170804
transform 1 0 17204 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _208_
timestamp 1693170804
transform -1 0 19136 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _209_
timestamp 1693170804
transform -1 0 17112 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _210_
timestamp 1693170804
transform -1 0 17388 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _211_
timestamp 1693170804
transform -1 0 19780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _212_
timestamp 1693170804
transform -1 0 16560 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_1  _213_
timestamp 1693170804
transform 1 0 17572 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_2  _214_
timestamp 1693170804
transform 1 0 17480 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _215_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _216_
timestamp 1693170804
transform 1 0 17112 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _217_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 17756 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _218_
timestamp 1693170804
transform 1 0 8372 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9752 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 13156 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1693170804
transform 1 0 13432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _223__2
timestamp 1693170804
transform 1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _224_
timestamp 1693170804
transform 1 0 3588 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1693170804
transform 1 0 5704 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _226_
timestamp 1693170804
transform -1 0 8924 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _227_
timestamp 1693170804
transform 1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228__3
timestamp 1693170804
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _229_
timestamp 1693170804
transform 1 0 3772 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1693170804
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _232_
timestamp 1693170804
transform 1 0 9016 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _233_
timestamp 1693170804
transform 1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234__4
timestamp 1693170804
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _235_
timestamp 1693170804
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _236_
timestamp 1693170804
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _237_
timestamp 1693170804
transform -1 0 12696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _241_
timestamp 1693170804
transform 1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _242_
timestamp 1693170804
transform 1 0 13156 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1693170804
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _244_
timestamp 1693170804
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _245_
timestamp 1693170804
transform 1 0 13156 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1693170804
transform -1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _247_
timestamp 1693170804
transform -1 0 3036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1693170804
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp 1693170804
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _250_
timestamp 1693170804
transform -1 0 2484 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1693170804
transform 1 0 1564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _252_
timestamp 1693170804
transform 1 0 3312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _253_
timestamp 1693170804
transform -1 0 3772 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1693170804
transform -1 0 3588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _255_
timestamp 1693170804
transform 1 0 1564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _256_
timestamp 1693170804
transform 1 0 6440 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1693170804
transform 1 0 6992 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _258_
timestamp 1693170804
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1693170804
transform 1 0 9752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _260_
timestamp 1693170804
transform -1 0 11408 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _261_
timestamp 1693170804
transform -1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _262_
timestamp 1693170804
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1693170804
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _264_
timestamp 1693170804
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _265_
timestamp 1693170804
transform 1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9660 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _267_
timestamp 1693170804
transform 1 0 9016 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 10396 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _269_
timestamp 1693170804
transform -1 0 9936 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _270_
timestamp 1693170804
transform -1 0 9660 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _271_
timestamp 1693170804
transform 1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _272_
timestamp 1693170804
transform 1 0 8740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 10396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 10120 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8372 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1693170804
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9108 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _278_
timestamp 1693170804
transform -1 0 10304 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10304 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _280_
timestamp 1693170804
transform 1 0 9384 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _281_
timestamp 1693170804
transform 1 0 9936 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _282_
timestamp 1693170804
transform 1 0 9660 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _283_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 10580 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9108 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _285_
timestamp 1693170804
transform -1 0 9384 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1693170804
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _287_
timestamp 1693170804
transform -1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1693170804
transform -1 0 12604 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _289_
timestamp 1693170804
transform -1 0 11408 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1693170804
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _291_
timestamp 1693170804
transform 1 0 11500 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _292_
timestamp 1693170804
transform 1 0 1380 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _293_
timestamp 1693170804
transform 1 0 3772 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _294_
timestamp 1693170804
transform -1 0 3680 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _295_
timestamp 1693170804
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _296_
timestamp 1693170804
transform 1 0 4876 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _297_
timestamp 1693170804
transform -1 0 5152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _298_
timestamp 1693170804
transform 1 0 5336 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _299_
timestamp 1693170804
transform -1 0 6440 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _300_
timestamp 1693170804
transform 1 0 6440 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _301_
timestamp 1693170804
transform -1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1693170804
transform 1 0 7176 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _303_
timestamp 1693170804
transform 1 0 7360 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _304_
timestamp 1693170804
transform 1 0 6900 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _305_
timestamp 1693170804
transform -1 0 8280 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _306_
timestamp 1693170804
transform -1 0 6256 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9844 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1693170804
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _309_
timestamp 1693170804
transform -1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _310_
timestamp 1693170804
transform -1 0 6256 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _311_
timestamp 1693170804
transform -1 0 5520 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _312_
timestamp 1693170804
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _313_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9660 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _314_
timestamp 1693170804
transform -1 0 9384 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1693170804
transform 1 0 8464 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _316_
timestamp 1693170804
transform 1 0 9108 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _317_
timestamp 1693170804
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _318__5
timestamp 1693170804
transform -1 0 12604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _319_
timestamp 1693170804
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _320_
timestamp 1693170804
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1693170804
transform 1 0 14444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _322_
timestamp 1693170804
transform 1 0 8464 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1693170804
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _324_
timestamp 1693170804
transform -1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _325__1
timestamp 1693170804
transform 1 0 4232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _326_
timestamp 1693170804
transform 1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1693170804
transform -1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1693170804
transform 1 0 4140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _329_
timestamp 1693170804
transform 1 0 8188 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _330_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _331_
timestamp 1693170804
transform 1 0 7820 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _332_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3772 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _333_
timestamp 1693170804
transform 1 0 2760 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _334_
timestamp 1693170804
transform -1 0 5060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4600 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _336_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _337_
timestamp 1693170804
transform 1 0 5336 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _338_
timestamp 1693170804
transform 1 0 6992 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _339_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 7820 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _340_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _341_
timestamp 1693170804
transform 1 0 7084 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _342_
timestamp 1693170804
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _345_
timestamp 1693170804
transform 1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _346_
timestamp 1693170804
transform 1 0 5520 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _347_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6440 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _348_
timestamp 1693170804
transform 1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _349_
timestamp 1693170804
transform -1 0 5244 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _350_
timestamp 1693170804
transform -1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _351_
timestamp 1693170804
transform 1 0 6348 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _352_
timestamp 1693170804
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _353_
timestamp 1693170804
transform 1 0 6900 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1693170804
transform -1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _355_
timestamp 1693170804
transform 1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _356_
timestamp 1693170804
transform -1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _357_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9108 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1693170804
transform -1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _359__6
timestamp 1693170804
transform -1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _360_
timestamp 1693170804
transform 1 0 4048 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  _361_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7728 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _362_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5612 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _363_
timestamp 1693170804
transform 1 0 6348 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _364_
timestamp 1693170804
transform 1 0 8924 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _365_
timestamp 1693170804
transform 1 0 6716 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _366_
timestamp 1693170804
transform -1 0 10396 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _367_
timestamp 1693170804
transform 1 0 9476 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _368_
timestamp 1693170804
transform 1 0 6992 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _369_
timestamp 1693170804
transform 1 0 7820 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _370_
timestamp 1693170804
transform 1 0 9292 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _371_
timestamp 1693170804
transform 1 0 9016 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _372_
timestamp 1693170804
transform 1 0 10304 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _373_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8004 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _374_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11500 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _375_
timestamp 1693170804
transform 1 0 9936 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _376_
timestamp 1693170804
transform 1 0 10212 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _377_
timestamp 1693170804
transform 1 0 14076 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _378_
timestamp 1693170804
transform 1 0 12236 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _379_
timestamp 1693170804
transform 1 0 11868 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _380_
timestamp 1693170804
transform 1 0 9476 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _381_
timestamp 1693170804
transform 1 0 14352 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _382_
timestamp 1693170804
transform 1 0 12512 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _383_
timestamp 1693170804
transform 1 0 14076 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _384_
timestamp 1693170804
transform 1 0 13064 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _385_
timestamp 1693170804
transform 1 0 14444 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _386_
timestamp 1693170804
transform 1 0 12604 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _387_
timestamp 1693170804
transform 1 0 9476 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _388_
timestamp 1693170804
transform -1 0 11040 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _389_
timestamp 1693170804
transform 1 0 3312 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _390_
timestamp 1693170804
transform -1 0 5796 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _391_
timestamp 1693170804
transform 1 0 1656 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _392_
timestamp 1693170804
transform 1 0 2760 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _393__21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _393_
timestamp 1693170804
transform 1 0 4324 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _394_
timestamp 1693170804
transform 1 0 5888 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _395_
timestamp 1693170804
transform 1 0 6808 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _396_
timestamp 1693170804
transform 1 0 2576 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _397_
timestamp 1693170804
transform 1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _398_
timestamp 1693170804
transform 1 0 1380 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _399_
timestamp 1693170804
transform 1 0 1840 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _400_
timestamp 1693170804
transform 1 0 1380 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _401_
timestamp 1693170804
transform 1 0 1840 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _402_
timestamp 1693170804
transform 1 0 3772 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _403_
timestamp 1693170804
transform -1 0 6072 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _404_
timestamp 1693170804
transform 1 0 1840 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _405_
timestamp 1693170804
transform 1 0 3772 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _406_
timestamp 1693170804
transform 1 0 5244 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _407_
timestamp 1693170804
transform 1 0 6716 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _408_
timestamp 1693170804
transform 1 0 2392 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _409_
timestamp 1693170804
transform 1 0 3772 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _410_
timestamp 1693170804
transform -1 0 8832 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _411_
timestamp 1693170804
transform 1 0 4508 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _412_
timestamp 1693170804
transform 1 0 8832 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _413_
timestamp 1693170804
transform 1 0 4508 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _414_
timestamp 1693170804
transform 1 0 6348 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _415_
timestamp 1693170804
transform 1 0 6348 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _416_
timestamp 1693170804
transform 1 0 6992 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 3312 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _418_
timestamp 1693170804
transform -1 0 3404 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _419_
timestamp 1693170804
transform -1 0 4324 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _420_
timestamp 1693170804
transform -1 0 5888 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _421_
timestamp 1693170804
transform 1 0 4692 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _422_
timestamp 1693170804
transform -1 0 7912 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _423_
timestamp 1693170804
transform 1 0 6256 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _424_
timestamp 1693170804
transform 1 0 10304 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _425_
timestamp 1693170804
transform 1 0 17572 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _426_
timestamp 1693170804
transform 1 0 18952 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _427_
timestamp 1693170804
transform 1 0 18952 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _428_
timestamp 1693170804
transform 1 0 18584 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _429_
timestamp 1693170804
transform 1 0 17572 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _430_
timestamp 1693170804
transform -1 0 18216 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _431_
timestamp 1693170804
transform 1 0 16652 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _432_
timestamp 1693170804
transform 1 0 15272 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _433_
timestamp 1693170804
transform 1 0 14260 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _434_
timestamp 1693170804
transform -1 0 15640 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _435_
timestamp 1693170804
transform -1 0 15640 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _436_
timestamp 1693170804
transform -1 0 13708 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _437_
timestamp 1693170804
transform -1 0 13616 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _438_
timestamp 1693170804
transform -1 0 18216 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _439_
timestamp 1693170804
transform 1 0 15640 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _440_
timestamp 1693170804
transform 1 0 14352 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _441_
timestamp 1693170804
transform -1 0 18216 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _442_
timestamp 1693170804
transform 1 0 14996 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _443_
timestamp 1693170804
transform 1 0 14168 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _444_
timestamp 1693170804
transform 1 0 14076 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _445_
timestamp 1693170804
transform 1 0 12880 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _446_
timestamp 1693170804
transform 1 0 11776 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _447_
timestamp 1693170804
transform -1 0 12880 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _448_
timestamp 1693170804
transform 1 0 11224 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _449_
timestamp 1693170804
transform 1 0 11132 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _450_
timestamp 1693170804
transform 1 0 9936 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _451_
timestamp 1693170804
transform -1 0 13064 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _452_
timestamp 1693170804
transform -1 0 13984 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _453_
timestamp 1693170804
transform 1 0 11592 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _454_
timestamp 1693170804
transform -1 0 13800 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _455_
timestamp 1693170804
transform 1 0 12144 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _456_
timestamp 1693170804
transform -1 0 13984 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _457_
timestamp 1693170804
transform 1 0 16744 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _458_
timestamp 1693170804
transform 1 0 18216 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _459_
timestamp 1693170804
transform 1 0 17388 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _460_
timestamp 1693170804
transform 1 0 18952 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _461_
timestamp 1693170804
transform 1 0 18492 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _462_
timestamp 1693170804
transform 1 0 17572 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _463_
timestamp 1693170804
transform 1 0 18584 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _464_
timestamp 1693170804
transform 1 0 17572 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _465_
timestamp 1693170804
transform 1 0 18216 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _466_
timestamp 1693170804
transform 1 0 16652 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _467_
timestamp 1693170804
transform 1 0 15916 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _468_
timestamp 1693170804
transform 1 0 15180 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _469_
timestamp 1693170804
transform -1 0 16192 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _470_
timestamp 1693170804
transform 1 0 15088 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _471_
timestamp 1693170804
transform -1 0 16560 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _472_
timestamp 1693170804
transform 1 0 14444 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _473_
timestamp 1693170804
transform -1 0 18492 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _474_
timestamp 1693170804
transform 1 0 18952 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _475_
timestamp 1693170804
transform 1 0 18584 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _476_
timestamp 1693170804
transform 1 0 18492 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _477_
timestamp 1693170804
transform 1 0 18584 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _478_
timestamp 1693170804
transform 1 0 18492 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _479_
timestamp 1693170804
transform 1 0 17572 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _480_
timestamp 1693170804
transform -1 0 19136 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _481_
timestamp 1693170804
transform 1 0 18216 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _482_
timestamp 1693170804
transform 1 0 16468 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _483_
timestamp 1693170804
transform -1 0 18216 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _484_
timestamp 1693170804
transform 1 0 15364 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _485_
timestamp 1693170804
transform -1 0 16192 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _486_
timestamp 1693170804
transform 1 0 15272 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _487_
timestamp 1693170804
transform -1 0 16192 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _488_
timestamp 1693170804
transform 1 0 13984 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 1693170804
transform 1 0 9016 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 1693170804
transform 1 0 10856 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 1693170804
transform 1 0 11408 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 1693170804
transform 1 0 13892 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 1693170804
transform 1 0 6992 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 1693170804
transform -1 0 10304 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 1693170804
transform 1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _496_
timestamp 1693170804
transform 1 0 6440 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__325__1_A
timestamp 1693170804
transform 1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__361__CLK
timestamp 1693170804
transform 1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__362__CLK
timestamp 1693170804
transform 1 0 5428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__363__CLK
timestamp 1693170804
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__364__CLK
timestamp 1693170804
transform 1 0 7912 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__365__CLK
timestamp 1693170804
transform 1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__366__CLK
timestamp 1693170804
transform -1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__367__CLK
timestamp 1693170804
transform 1 0 10120 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__368__CLK
timestamp 1693170804
transform 1 0 6808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__369__CLK
timestamp 1693170804
transform 1 0 7636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__370__CLK
timestamp 1693170804
transform 1 0 8188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__371__CLK
timestamp 1693170804
transform 1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__372__CLK
timestamp 1693170804
transform -1 0 10580 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__373__CLK
timestamp 1693170804
transform 1 0 7820 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__396__CLK
timestamp 1693170804
transform 1 0 2392 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__CLK
timestamp 1693170804
transform 1 0 3588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__CLK
timestamp 1693170804
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__406__CLK
timestamp 1693170804
transform 1 0 5060 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__407__CLK
timestamp 1693170804
transform 1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__408__CLK
timestamp 1693170804
transform 1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__409__CLK
timestamp 1693170804
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__410__CLK
timestamp 1693170804
transform 1 0 6808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__411__CLK
timestamp 1693170804
transform 1 0 4324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__412__CLK
timestamp 1693170804
transform 1 0 8004 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__417__CLK
timestamp 1693170804
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__418__CLK
timestamp 1693170804
transform 1 0 3128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__419__CLK
timestamp 1693170804
transform -1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__420__CLK
timestamp 1693170804
transform 1 0 4140 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__CLK
timestamp 1693170804
transform 1 0 4508 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__CLK
timestamp 1693170804
transform 1 0 5888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__CLK
timestamp 1693170804
transform -1 0 5980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__CLK
timestamp 1693170804
transform -1 0 10304 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__026_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11316 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__041_
timestamp 1693170804
transform 1 0 6348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__045_
timestamp 1693170804
transform 1 0 9016 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLKMUX.clko
timestamp 1693170804
transform 1 0 12052 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLKMUX.clko1
timestamp 1693170804
transform -1 0 13156 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_PoR.clk_div\[8\]
timestamp 1693170804
transform 1 0 14536 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__026_
timestamp 1693170804
transform -1 0 10764 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__041_
timestamp 1693170804
transform -1 0 4600 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__045_
timestamp 1693170804
transform -1 0 8832 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CLKMUX.clko
timestamp 1693170804
transform -1 0 10764 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CLKMUX.clko1
timestamp 1693170804
transform -1 0 10028 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__026_
timestamp 1693170804
transform 1 0 10856 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__041_
timestamp 1693170804
transform 1 0 5152 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__045_
timestamp 1693170804
transform -1 0 10028 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CLKMUX.clko
timestamp 1693170804
transform 1 0 14076 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CLKMUX.clko1
timestamp 1693170804
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_PoR.clk_div\[8\]
timestamp 1693170804
transform -1 0 15916 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_PoR.clk_div\[8\]
timestamp 1693170804
transform 1 0 13616 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_PoR.clk_div\[8\]
timestamp 1693170804
transform 1 0 16652 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_PoR.clk_div\[8\]
timestamp 1693170804
transform 1 0 16284 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_PoR.clk_div\[8\]
timestamp 1693170804
transform -1 0 13340 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_PoR.clk_div\[8\]
timestamp 1693170804
transform -1 0 13340 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_PoR.clk_div\[8\]
timestamp 1693170804
transform 1 0 16652 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_PoR.clk_div\[8\]
timestamp 1693170804
transform 1 0 16652 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12144 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1693170804
transform -1 0 6900 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1693170804
transform -1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1693170804
transform -1 0 7728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1693170804
transform -1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1693170804
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1693170804
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 1693170804
transform -1 0 12052 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1693170804
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1693170804
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6348 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_63
timestamp 1693170804
transform 1 0 6900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_125
timestamp 1693170804
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_134
timestamp 1693170804
transform 1 0 13432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1693170804
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1693170804
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153
timestamp 1693170804
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_161
timestamp 1693170804
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1693170804
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1693170804
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1693170804
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1693170804
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_209
timestamp 1693170804
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1693170804
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_15
timestamp 1693170804
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_23
timestamp 1693170804
transform 1 0 3220 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_44
timestamp 1693170804
transform 1 0 5152 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1693170804
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_69
timestamp 1693170804
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_77
timestamp 1693170804
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_100
timestamp 1693170804
transform 1 0 10304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1693170804
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_164
timestamp 1693170804
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1693170804
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1693170804
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1693170804
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_205
timestamp 1693170804
transform 1 0 19964 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1693170804
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1693170804
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1693170804
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1693170804
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_51
timestamp 1693170804
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_63
timestamp 1693170804
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1693170804
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_98
timestamp 1693170804
transform 1 0 10120 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_115
timestamp 1693170804
transform 1 0 11684 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_161
timestamp 1693170804
transform 1 0 15916 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_173
timestamp 1693170804
transform 1 0 17020 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_185
timestamp 1693170804
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_193
timestamp 1693170804
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1693170804
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_209
timestamp 1693170804
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1693170804
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1693170804
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_27
timestamp 1693170804
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_34
timestamp 1693170804
transform 1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_46
timestamp 1693170804
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1693170804
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1693170804
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1693170804
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_94
timestamp 1693170804
transform 1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_129
timestamp 1693170804
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_150
timestamp 1693170804
transform 1 0 14904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_162
timestamp 1693170804
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1693170804
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1693170804
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1693170804
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_205
timestamp 1693170804
transform 1 0 19964 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1693170804
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1693170804
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1693170804
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_29
timestamp 1693170804
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_39
timestamp 1693170804
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_43
timestamp 1693170804
transform 1 0 5060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_48
timestamp 1693170804
transform 1 0 5520 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_59
timestamp 1693170804
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_71
timestamp 1693170804
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1693170804
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1693170804
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_126
timestamp 1693170804
transform 1 0 12696 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_132
timestamp 1693170804
transform 1 0 13248 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1693170804
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1693170804
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1693170804
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1693170804
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1693170804
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1693170804
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1693170804
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1693170804
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_209
timestamp 1693170804
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_3
timestamp 1693170804
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_27
timestamp 1693170804
transform 1 0 3588 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1693170804
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_79
timestamp 1693170804
transform 1 0 8372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1693170804
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_148
timestamp 1693170804
transform 1 0 14720 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_160
timestamp 1693170804
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1693170804
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1693170804
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1693170804
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_205
timestamp 1693170804
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1693170804
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1693170804
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 1693170804
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_72
timestamp 1693170804
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_178
timestamp 1693170804
transform 1 0 17480 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_190
timestamp 1693170804
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1693170804
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_209
timestamp 1693170804
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1693170804
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_38
timestamp 1693170804
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_50
timestamp 1693170804
transform 1 0 5704 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_100
timestamp 1693170804
transform 1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_106
timestamp 1693170804
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_121
timestamp 1693170804
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_165
timestamp 1693170804
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_203
timestamp 1693170804
transform 1 0 19780 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1693170804
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1693170804
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1693170804
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_29
timestamp 1693170804
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_72
timestamp 1693170804
transform 1 0 7728 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_105
timestamp 1693170804
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_110
timestamp 1693170804
transform 1 0 11224 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_122
timestamp 1693170804
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_134
timestamp 1693170804
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1693170804
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_177
timestamp 1693170804
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1693170804
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_209
timestamp 1693170804
transform 1 0 20332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1693170804
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_11
timestamp 1693170804
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_34
timestamp 1693170804
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_48
timestamp 1693170804
transform 1 0 5520 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_65
timestamp 1693170804
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_97
timestamp 1693170804
transform 1 0 10028 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1693170804
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_137
timestamp 1693170804
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_145
timestamp 1693170804
transform 1 0 14444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_164
timestamp 1693170804
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1693170804
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_176
timestamp 1693170804
transform 1 0 17296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_188
timestamp 1693170804
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_207
timestamp 1693170804
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_16
timestamp 1693170804
transform 1 0 2576 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_24
timestamp 1693170804
transform 1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_49
timestamp 1693170804
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1693170804
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 1693170804
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_149
timestamp 1693170804
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_210
timestamp 1693170804
transform 1 0 20424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1693170804
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1693170804
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_27
timestamp 1693170804
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_45
timestamp 1693170804
transform 1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1693170804
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_71
timestamp 1693170804
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_161
timestamp 1693170804
transform 1 0 15916 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1693170804
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_206
timestamp 1693170804
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_210
timestamp 1693170804
transform 1 0 20424 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 1693170804
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_13
timestamp 1693170804
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1693170804
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1693170804
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1693170804
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_44
timestamp 1693170804
transform 1 0 5152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_51
timestamp 1693170804
transform 1 0 5796 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_59
timestamp 1693170804
transform 1 0 6532 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_64
timestamp 1693170804
transform 1 0 6992 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_76
timestamp 1693170804
transform 1 0 8096 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1693170804
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_89
timestamp 1693170804
transform 1 0 9292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_137
timestamp 1693170804
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_141
timestamp 1693170804
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_149
timestamp 1693170804
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_168
timestamp 1693170804
transform 1 0 16560 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_176
timestamp 1693170804
transform 1 0 17296 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1693170804
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1693170804
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1693170804
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_209
timestamp 1693170804
transform 1 0 20332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_3
timestamp 1693170804
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_11
timestamp 1693170804
transform 1 0 2116 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_17
timestamp 1693170804
transform 1 0 2668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_21
timestamp 1693170804
transform 1 0 3036 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_25
timestamp 1693170804
transform 1 0 3404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_46
timestamp 1693170804
transform 1 0 5336 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1693170804
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_76
timestamp 1693170804
transform 1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_94
timestamp 1693170804
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_104
timestamp 1693170804
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp 1693170804
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_119
timestamp 1693170804
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_126
timestamp 1693170804
transform 1 0 12696 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_138
timestamp 1693170804
transform 1 0 13800 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_144
timestamp 1693170804
transform 1 0 14352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_162
timestamp 1693170804
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_169
timestamp 1693170804
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1693170804
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_7
timestamp 1693170804
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_57
timestamp 1693170804
transform 1 0 6348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1693170804
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_90
timestamp 1693170804
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_97
timestamp 1693170804
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_101
timestamp 1693170804
transform 1 0 10396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_105
timestamp 1693170804
transform 1 0 10764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_141
timestamp 1693170804
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_161
timestamp 1693170804
transform 1 0 15916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_169
timestamp 1693170804
transform 1 0 16652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_197
timestamp 1693170804
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_205
timestamp 1693170804
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1693170804
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_13
timestamp 1693170804
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_17
timestamp 1693170804
transform 1 0 2668 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_38
timestamp 1693170804
transform 1 0 4600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_102
timestamp 1693170804
transform 1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_117
timestamp 1693170804
transform 1 0 11868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_159
timestamp 1693170804
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1693170804
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_210
timestamp 1693170804
transform 1 0 20424 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_6
timestamp 1693170804
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 1693170804
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1693170804
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1693170804
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_41
timestamp 1693170804
transform 1 0 4876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_65
timestamp 1693170804
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_69
timestamp 1693170804
transform 1 0 7452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_72
timestamp 1693170804
transform 1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1693170804
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1693170804
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_161
timestamp 1693170804
transform 1 0 15916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_190
timestamp 1693170804
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_203
timestamp 1693170804
transform 1 0 19780 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_23
timestamp 1693170804
transform 1 0 3220 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_29
timestamp 1693170804
transform 1 0 3772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_41
timestamp 1693170804
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1693170804
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1693170804
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_69
timestamp 1693170804
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_77
timestamp 1693170804
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_83
timestamp 1693170804
transform 1 0 8740 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_91
timestamp 1693170804
transform 1 0 9476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_97
timestamp 1693170804
transform 1 0 10028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_105
timestamp 1693170804
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1693170804
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 1693170804
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_156
timestamp 1693170804
transform 1 0 15456 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1693170804
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_179
timestamp 1693170804
transform 1 0 17572 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_191
timestamp 1693170804
transform 1 0 18676 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1693170804
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_37
timestamp 1693170804
transform 1 0 4508 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_49
timestamp 1693170804
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_61
timestamp 1693170804
transform 1 0 6716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_73
timestamp 1693170804
transform 1 0 7820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1693170804
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_93
timestamp 1693170804
transform 1 0 9660 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_105
timestamp 1693170804
transform 1 0 10764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_117
timestamp 1693170804
transform 1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_125
timestamp 1693170804
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_134
timestamp 1693170804
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_175
timestamp 1693170804
transform 1 0 17204 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_208
timestamp 1693170804
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_3
timestamp 1693170804
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_15
timestamp 1693170804
transform 1 0 2484 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_66
timestamp 1693170804
transform 1 0 7176 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_72
timestamp 1693170804
transform 1 0 7728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_103
timestamp 1693170804
transform 1 0 10580 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_119
timestamp 1693170804
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_137
timestamp 1693170804
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_164
timestamp 1693170804
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_186
timestamp 1693170804
transform 1 0 18216 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_3
timestamp 1693170804
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_11
timestamp 1693170804
transform 1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_16
timestamp 1693170804
transform 1 0 2576 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1693170804
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp 1693170804
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1693170804
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1693170804
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_90
timestamp 1693170804
transform 1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_131
timestamp 1693170804
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1693170804
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_160
timestamp 1693170804
transform 1 0 15824 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_168
timestamp 1693170804
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_186
timestamp 1693170804
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1693170804
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1693170804
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_209
timestamp 1693170804
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1693170804
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_15
timestamp 1693170804
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_49
timestamp 1693170804
transform 1 0 5612 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_85
timestamp 1693170804
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_89
timestamp 1693170804
transform 1 0 9292 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_99
timestamp 1693170804
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_103
timestamp 1693170804
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1693170804
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_133
timestamp 1693170804
transform 1 0 13340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_145
timestamp 1693170804
transform 1 0 14444 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1693170804
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 1693170804
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_207
timestamp 1693170804
transform 1 0 20148 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_3
timestamp 1693170804
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1693170804
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_41
timestamp 1693170804
transform 1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1693170804
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_106
timestamp 1693170804
transform 1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_110
timestamp 1693170804
transform 1 0 11224 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_128
timestamp 1693170804
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1693170804
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_153
timestamp 1693170804
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_177
timestamp 1693170804
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1693170804
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_209
timestamp 1693170804
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_23
timestamp 1693170804
transform 1 0 3220 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1693170804
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_77
timestamp 1693170804
transform 1 0 8188 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_83
timestamp 1693170804
transform 1 0 8740 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_86
timestamp 1693170804
transform 1 0 9016 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_92
timestamp 1693170804
transform 1 0 9568 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 1693170804
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1693170804
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_113
timestamp 1693170804
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_133
timestamp 1693170804
transform 1 0 13340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_141
timestamp 1693170804
transform 1 0 14076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_159
timestamp 1693170804
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1693170804
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1693170804
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 1693170804
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_206
timestamp 1693170804
transform 1 0 20056 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_210
timestamp 1693170804
transform 1 0 20424 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 1693170804
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_7
timestamp 1693170804
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_11
timestamp 1693170804
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_23
timestamp 1693170804
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1693170804
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_29
timestamp 1693170804
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_36
timestamp 1693170804
transform 1 0 4416 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_48
timestamp 1693170804
transform 1 0 5520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_56
timestamp 1693170804
transform 1 0 6256 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_67
timestamp 1693170804
transform 1 0 7268 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1693170804
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1693170804
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1693170804
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1693170804
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_109
timestamp 1693170804
transform 1 0 11132 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_165
timestamp 1693170804
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_173
timestamp 1693170804
transform 1 0 17020 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_191
timestamp 1693170804
transform 1 0 18676 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1693170804
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1693170804
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_209
timestamp 1693170804
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_18
timestamp 1693170804
transform 1 0 2760 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_28
timestamp 1693170804
transform 1 0 3680 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_32
timestamp 1693170804
transform 1 0 4048 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_35
timestamp 1693170804
transform 1 0 4324 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_44
timestamp 1693170804
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1693170804
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_69
timestamp 1693170804
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_101
timestamp 1693170804
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1693170804
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1693170804
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_125
timestamp 1693170804
transform 1 0 12604 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_186
timestamp 1693170804
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_207
timestamp 1693170804
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_7
timestamp 1693170804
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_25
timestamp 1693170804
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_34
timestamp 1693170804
transform 1 0 4232 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_73
timestamp 1693170804
transform 1 0 7820 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_88
timestamp 1693170804
transform 1 0 9200 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_126
timestamp 1693170804
transform 1 0 12696 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1693170804
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_141
timestamp 1693170804
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_149
timestamp 1693170804
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_164
timestamp 1693170804
transform 1 0 16192 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_176
timestamp 1693170804
transform 1 0 17296 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_187
timestamp 1693170804
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_204
timestamp 1693170804
transform 1 0 19872 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_210
timestamp 1693170804
transform 1 0 20424 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_3
timestamp 1693170804
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1693170804
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_61
timestamp 1693170804
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_83
timestamp 1693170804
transform 1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_94
timestamp 1693170804
transform 1 0 9752 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_98
timestamp 1693170804
transform 1 0 10120 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_107
timestamp 1693170804
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1693170804
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1693170804
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_131
timestamp 1693170804
transform 1 0 13156 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_142
timestamp 1693170804
transform 1 0 14168 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_154
timestamp 1693170804
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1693170804
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_169
timestamp 1693170804
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_189
timestamp 1693170804
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_193
timestamp 1693170804
transform 1 0 18860 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_3
timestamp 1693170804
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_24
timestamp 1693170804
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_40
timestamp 1693170804
transform 1 0 4784 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_52
timestamp 1693170804
transform 1 0 5888 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_64
timestamp 1693170804
transform 1 0 6992 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_76
timestamp 1693170804
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1693170804
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_93
timestamp 1693170804
transform 1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1693170804
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_141
timestamp 1693170804
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_164
timestamp 1693170804
transform 1 0 16192 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_176
timestamp 1693170804
transform 1 0 17296 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_184
timestamp 1693170804
transform 1 0 18032 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_203
timestamp 1693170804
transform 1 0 19780 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_3
timestamp 1693170804
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_9
timestamp 1693170804
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_14
timestamp 1693170804
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_26
timestamp 1693170804
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_38
timestamp 1693170804
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_50
timestamp 1693170804
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_57
timestamp 1693170804
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_61
timestamp 1693170804
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_64
timestamp 1693170804
transform 1 0 6992 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_76
timestamp 1693170804
transform 1 0 8096 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_82
timestamp 1693170804
transform 1 0 8648 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_96
timestamp 1693170804
transform 1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_100
timestamp 1693170804
transform 1 0 10304 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 1693170804
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_121
timestamp 1693170804
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_157
timestamp 1693170804
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1693170804
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_174
timestamp 1693170804
transform 1 0 17112 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_185
timestamp 1693170804
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_189
timestamp 1693170804
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_207
timestamp 1693170804
transform 1 0 20148 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_3
timestamp 1693170804
transform 1 0 1380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_9
timestamp 1693170804
transform 1 0 1932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_22
timestamp 1693170804
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1693170804
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_41
timestamp 1693170804
transform 1 0 4876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_63
timestamp 1693170804
transform 1 0 6900 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 1693170804
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_111
timestamp 1693170804
transform 1 0 11316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_131
timestamp 1693170804
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1693170804
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1693170804
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_153
timestamp 1693170804
transform 1 0 15180 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_177
timestamp 1693170804
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 1693170804
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp 1693170804
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_209
timestamp 1693170804
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1693170804
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_35
timestamp 1693170804
transform 1 0 4324 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_74
timestamp 1693170804
transform 1 0 7912 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_101
timestamp 1693170804
transform 1 0 10396 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp 1693170804
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_138
timestamp 1693170804
transform 1 0 13800 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_150
timestamp 1693170804
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_162
timestamp 1693170804
transform 1 0 16008 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_206
timestamp 1693170804
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_210
timestamp 1693170804
transform 1 0 20424 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1693170804
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1693170804
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1693170804
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_33
timestamp 1693170804
transform 1 0 4140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_45
timestamp 1693170804
transform 1 0 5244 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_51
timestamp 1693170804
transform 1 0 5796 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_69
timestamp 1693170804
transform 1 0 7452 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_77
timestamp 1693170804
transform 1 0 8188 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1693170804
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_100
timestamp 1693170804
transform 1 0 10304 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_112
timestamp 1693170804
transform 1 0 11408 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_137
timestamp 1693170804
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_146
timestamp 1693170804
transform 1 0 14536 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_154
timestamp 1693170804
transform 1 0 15272 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1693170804
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_209
timestamp 1693170804
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1693170804
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1693170804
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_27
timestamp 1693170804
transform 1 0 3588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_38
timestamp 1693170804
transform 1 0 4600 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_50
timestamp 1693170804
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1693170804
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_101
timestamp 1693170804
transform 1 0 10396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1693170804
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1693170804
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_138
timestamp 1693170804
transform 1 0 13800 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_146
timestamp 1693170804
transform 1 0 14536 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_164
timestamp 1693170804
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_203
timestamp 1693170804
transform 1 0 19780 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1693170804
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1693170804
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1693170804
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_29
timestamp 1693170804
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_35
timestamp 1693170804
transform 1 0 4324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_40
timestamp 1693170804
transform 1 0 4784 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_48
timestamp 1693170804
transform 1 0 5520 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_78
timestamp 1693170804
transform 1 0 8280 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1693170804
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_85
timestamp 1693170804
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_89
timestamp 1693170804
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_93
timestamp 1693170804
transform 1 0 9660 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_97
timestamp 1693170804
transform 1 0 10028 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_117
timestamp 1693170804
transform 1 0 11868 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1693170804
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1693170804
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_165
timestamp 1693170804
transform 1 0 16284 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_184
timestamp 1693170804
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1693170804
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_209
timestamp 1693170804
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1693170804
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1693170804
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_27
timestamp 1693170804
transform 1 0 3588 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1693170804
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1693170804
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1693170804
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_57
timestamp 1693170804
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_71
timestamp 1693170804
transform 1 0 7636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_83
timestamp 1693170804
transform 1 0 8740 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_85
timestamp 1693170804
transform 1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_93
timestamp 1693170804
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_108
timestamp 1693170804
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1693170804
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1693170804
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_137
timestamp 1693170804
transform 1 0 13708 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_145
timestamp 1693170804
transform 1 0 14444 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_157
timestamp 1693170804
transform 1 0 15548 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_165
timestamp 1693170804
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1693170804
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_181
timestamp 1693170804
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_189
timestamp 1693170804
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_195
timestamp 1693170804
transform 1 0 19044 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_197
timestamp 1693170804
transform 1 0 19228 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_205
timestamp 1693170804
transform 1 0 19964 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 13432 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold2
timestamp 1693170804
transform -1 0 12420 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1693170804
transform -1 0 11500 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1693170804
transform -1 0 13984 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1693170804
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1693170804
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1693170804
transform -1 0 7728 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1693170804
transform -1 0 9108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1693170804
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1693170804
transform -1 0 14076 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1693170804
transform -1 0 5796 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1693170804
transform 1 0 2024 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1693170804
transform 1 0 6440 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold14
timestamp 1693170804
transform -1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1693170804
transform 1 0 2024 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1693170804
transform -1 0 11408 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1693170804
transform -1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1693170804
transform -1 0 10948 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1693170804
transform -1 0 12512 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1693170804
transform -1 0 12236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1693170804
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1693170804
transform -1 0 10028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1693170804
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1693170804
transform -1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1693170804
transform -1 0 11224 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1693170804
transform -1 0 6348 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1693170804
transform -1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1693170804
transform -1 0 13432 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1693170804
transform 1 0 14076 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1693170804
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1693170804
transform -1 0 20516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1693170804
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1693170804
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1693170804
transform -1 0 19044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1693170804
transform 1 0 10396 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1693170804
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1693170804
transform 1 0 3772 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1693170804
transform -1 0 20516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1693170804
transform 1 0 20148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1693170804
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_36
timestamp 1693170804
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_37
timestamp 1693170804
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_38
timestamp 1693170804
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_39
timestamp 1693170804
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_40
timestamp 1693170804
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 20792 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_41
timestamp 1693170804
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_42
timestamp 1693170804
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 20792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_43
timestamp 1693170804
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_44
timestamp 1693170804
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 20792 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_45
timestamp 1693170804
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_46
timestamp 1693170804
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_47
timestamp 1693170804
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1693170804
transform -1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_48
timestamp 1693170804
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1693170804
transform -1 0 20792 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_49
timestamp 1693170804
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1693170804
transform -1 0 20792 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_50
timestamp 1693170804
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1693170804
transform -1 0 20792 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_51
timestamp 1693170804
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1693170804
transform -1 0 20792 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_52
timestamp 1693170804
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1693170804
transform -1 0 20792 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_53
timestamp 1693170804
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1693170804
transform -1 0 20792 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_54
timestamp 1693170804
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1693170804
transform -1 0 20792 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_55
timestamp 1693170804
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1693170804
transform -1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_56
timestamp 1693170804
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1693170804
transform -1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_57
timestamp 1693170804
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1693170804
transform -1 0 20792 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_58
timestamp 1693170804
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1693170804
transform -1 0 20792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_59
timestamp 1693170804
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1693170804
transform -1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_60
timestamp 1693170804
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1693170804
transform -1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_61
timestamp 1693170804
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1693170804
transform -1 0 20792 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_62
timestamp 1693170804
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1693170804
transform -1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_63
timestamp 1693170804
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1693170804
transform -1 0 20792 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_64
timestamp 1693170804
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1693170804
transform -1 0 20792 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_65
timestamp 1693170804
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1693170804
transform -1 0 20792 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_66
timestamp 1693170804
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1693170804
transform -1 0 20792 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_67
timestamp 1693170804
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1693170804
transform -1 0 20792 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_68
timestamp 1693170804
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1693170804
transform -1 0 20792 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_69
timestamp 1693170804
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1693170804
transform -1 0 20792 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_70
timestamp 1693170804
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1693170804
transform -1 0 20792 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_71
timestamp 1693170804
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1693170804
transform -1 0 20792 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  PoR.ROSC_CLKBUF_0
timestamp 1693170804
transform -1 0 2484 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  PoR.ROSC_CLKBUF_1
timestamp 1693170804
transform 1 0 1472 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYBUF_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_0.clkdlybuf
timestamp 1693170804
transform -1 0 4600 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_0.clkinv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 4784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_1.clkdlybuf
timestamp 1693170804
transform 1 0 3220 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_1.clkinv
timestamp 1693170804
transform -1 0 4140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_2.clkdlybuf
timestamp 1693170804
transform -1 0 3220 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_2.clkinv
timestamp 1693170804
transform 1 0 3956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_3.clkdlybuf
timestamp 1693170804
transform -1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_3.clkinv
timestamp 1693170804
transform 1 0 2760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_4.clkdlybuf
timestamp 1693170804
transform -1 0 2300 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_4.clkinv
timestamp 1693170804
transform -1 0 2392 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  PoR.ROSC_DLYINV_5.clkdlybuf
timestamp 1693170804
transform 1 0 1564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  PoR.ROSC_DLYINV_5.clkinv
timestamp 1693170804
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  PoR.ROSC_DLYINV_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform -1 0 2576 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1693170804
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1693170804
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 1693170804
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 1693170804
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 1693170804
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 1693170804
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 1693170804
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 1693170804
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 1693170804
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_82
timestamp 1693170804
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_83
timestamp 1693170804
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 1693170804
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 1693170804
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_86
timestamp 1693170804
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_87
timestamp 1693170804
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_88
timestamp 1693170804
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_89
timestamp 1693170804
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_90
timestamp 1693170804
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_91
timestamp 1693170804
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_92
timestamp 1693170804
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_93
timestamp 1693170804
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_94
timestamp 1693170804
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_95
timestamp 1693170804
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_96
timestamp 1693170804
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_97
timestamp 1693170804
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_98
timestamp 1693170804
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_99
timestamp 1693170804
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_100
timestamp 1693170804
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_101
timestamp 1693170804
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp 1693170804
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_103
timestamp 1693170804
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_104
timestamp 1693170804
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_105
timestamp 1693170804
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_106
timestamp 1693170804
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_107
timestamp 1693170804
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_108
timestamp 1693170804
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp 1693170804
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_110
timestamp 1693170804
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_111
timestamp 1693170804
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_112
timestamp 1693170804
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp 1693170804
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_114
timestamp 1693170804
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_115
timestamp 1693170804
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_116
timestamp 1693170804
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_117
timestamp 1693170804
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_118
timestamp 1693170804
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_119
timestamp 1693170804
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_120
timestamp 1693170804
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_121
timestamp 1693170804
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_122
timestamp 1693170804
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_123
timestamp 1693170804
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_124
timestamp 1693170804
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_125
timestamp 1693170804
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_126
timestamp 1693170804
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_127
timestamp 1693170804
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_128
timestamp 1693170804
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_129
timestamp 1693170804
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_130
timestamp 1693170804
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_131
timestamp 1693170804
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_132
timestamp 1693170804
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_133
timestamp 1693170804
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_134
timestamp 1693170804
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_135
timestamp 1693170804
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_136
timestamp 1693170804
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_137
timestamp 1693170804
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_138
timestamp 1693170804
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_139
timestamp 1693170804
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_140
timestamp 1693170804
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_141
timestamp 1693170804
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_142
timestamp 1693170804
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_143
timestamp 1693170804
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_144
timestamp 1693170804
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_145
timestamp 1693170804
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_146
timestamp 1693170804
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_147
timestamp 1693170804
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_148
timestamp 1693170804
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_149
timestamp 1693170804
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_150
timestamp 1693170804
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_151
timestamp 1693170804
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_152
timestamp 1693170804
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_153
timestamp 1693170804
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_154
timestamp 1693170804
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_155
timestamp 1693170804
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_156
timestamp 1693170804
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_157
timestamp 1693170804
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_158
timestamp 1693170804
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_159
timestamp 1693170804
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_160
timestamp 1693170804
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_161
timestamp 1693170804
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_162
timestamp 1693170804
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_163
timestamp 1693170804
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_164
timestamp 1693170804
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_165
timestamp 1693170804
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_166
timestamp 1693170804
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_167
timestamp 1693170804
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_168
timestamp 1693170804
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_169
timestamp 1693170804
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_170
timestamp 1693170804
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_171
timestamp 1693170804
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_172
timestamp 1693170804
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_173
timestamp 1693170804
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_174
timestamp 1693170804
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_175
timestamp 1693170804
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_176
timestamp 1693170804
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_177
timestamp 1693170804
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_178
timestamp 1693170804
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_179
timestamp 1693170804
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_180
timestamp 1693170804
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_181
timestamp 1693170804
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_182
timestamp 1693170804
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_183
timestamp 1693170804
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_184
timestamp 1693170804
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_185
timestamp 1693170804
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_186
timestamp 1693170804
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_187
timestamp 1693170804
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_188
timestamp 1693170804
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_189
timestamp 1693170804
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_190
timestamp 1693170804
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1693170804
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1693170804
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1693170804
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_194
timestamp 1693170804
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_195
timestamp 1693170804
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_196
timestamp 1693170804
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_197
timestamp 1693170804
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_198
timestamp 1693170804
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_199
timestamp 1693170804
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_200
timestamp 1693170804
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_201
timestamp 1693170804
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_202
timestamp 1693170804
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_203
timestamp 1693170804
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_204
timestamp 1693170804
transform 1 0 19136 0 -1 21760
box -38 -48 130 592
<< labels >>
flabel metal3 s 21146 15648 21946 15768 0 FreeSans 480 0 0 0 clk
port 0 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 clk_div[0]
port 1 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 clk_div[1]
port 2 nsew signal input
flabel metal2 s 13542 23290 13598 24090 0 FreeSans 224 90 0 0 one
port 3 nsew signal input
flabel metal2 s 8390 23290 8446 24090 0 FreeSans 224 90 0 0 por_fb_in
port 4 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 por_fb_out
port 5 nsew signal tristate
flabel metal3 s 21146 21088 21946 21208 0 FreeSans 480 0 0 0 por_n
port 6 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 rst_n
port 7 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 sel_mux0
port 8 nsew signal input
flabel metal3 s 21146 4768 21946 4888 0 FreeSans 480 0 0 0 sel_mux1
port 9 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 sel_mux2
port 10 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 sel_rosc[0]
port 11 nsew signal input
flabel metal2 s 18694 23290 18750 24090 0 FreeSans 224 90 0 0 sel_rosc[1]
port 12 nsew signal input
flabel metal4 s 4208 2128 4528 21808 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 10208 2128 10528 21808 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 16208 2128 16528 21808 0 FreeSans 1920 90 0 0 vccd1
port 13 nsew power bidirectional
flabel metal4 s 7208 2128 7528 21808 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal4 s 13208 2128 13528 21808 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal4 s 19208 2128 19528 21808 0 FreeSans 1920 90 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 xclk0
port 15 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 xclk1
port 16 nsew signal input
flabel metal2 s 3238 23290 3294 24090 0 FreeSans 224 90 0 0 xrst_n
port 17 nsew signal input
flabel metal3 s 21146 10208 21946 10328 0 FreeSans 480 0 0 0 zero
port 18 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 21946 24090
<< end >>
